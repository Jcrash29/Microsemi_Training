`timescale 1 ns/100 ps
// Version: v11.7 SP1 11.7.1.11


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module MSS_025(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MGPIO25A_IN,
       MGPIO26A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_CTS_MGPIO13B_IN,
       MMUART1_DCD_MGPIO16B_IN,
       MMUART1_DSR_MGPIO14B_IN,
       MMUART1_DTR_MGPIO12B_IN,
       MMUART1_RI_MGPIO15B_IN,
       MMUART1_RTS_MGPIO11B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI0_SS4_MGPIO19A_IN,
       SPI0_SS5_MGPIO20A_IN,
       SPI0_SS6_MGPIO21A_IN,
       SPI0_SS7_MGPIO22A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MGPIO25A_OUT,
       MGPIO26A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_CTS_MGPIO13B_OUT,
       MMUART1_DCD_MGPIO16B_OUT,
       MMUART1_DSR_MGPIO14B_OUT,
       MMUART1_DTR_MGPIO12B_OUT,
       MMUART1_RI_MGPIO15B_OUT,
       MMUART1_RTS_MGPIO11B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI0_SS4_MGPIO19A_OUT,
       SPI0_SS5_MGPIO20A_OUT,
       SPI0_SS6_MGPIO21A_OUT,
       SPI0_SS7_MGPIO22A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MGPIO25A_OE,
       MGPIO26A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_CTS_MGPIO13B_OE,
       MMUART1_DCD_MGPIO16B_OE,
       MMUART1_DSR_MGPIO14B_OE,
       MMUART1_DTR_MGPIO12B_OE,
       MMUART1_RI_MGPIO15B_OE,
       MMUART1_RTS_MGPIO11B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI0_SS4_MGPIO19A_OE,
       SPI0_SS5_MGPIO20A_OE,
       SPI0_SS6_MGPIO21A_OE,
       SPI0_SS7_MGPIO22A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MGPIO25A_IN;
input  MGPIO26A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_CTS_MGPIO13B_IN;
input  MMUART1_DCD_MGPIO16B_IN;
input  MMUART1_DSR_MGPIO14B_IN;
input  MMUART1_DTR_MGPIO12B_IN;
input  MMUART1_RI_MGPIO15B_IN;
input  MMUART1_RTS_MGPIO11B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI0_SS4_MGPIO19A_IN;
input  SPI0_SS5_MGPIO20A_IN;
input  SPI0_SS6_MGPIO21A_IN;
input  SPI0_SS7_MGPIO22A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MGPIO25A_OUT;
output MGPIO26A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_CTS_MGPIO13B_OUT;
output MMUART1_DCD_MGPIO16B_OUT;
output MMUART1_DSR_MGPIO14B_OUT;
output MMUART1_DTR_MGPIO12B_OUT;
output MMUART1_RI_MGPIO15B_OUT;
output MMUART1_RTS_MGPIO11B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI0_SS4_MGPIO19A_OUT;
output SPI0_SS5_MGPIO20A_OUT;
output SPI0_SS6_MGPIO21A_OUT;
output SPI0_SS7_MGPIO22A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MGPIO25A_OE;
output MGPIO26A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_CTS_MGPIO13B_OE;
output MMUART1_DCD_MGPIO16B_OE;
output MMUART1_DSR_MGPIO14B_OE;
output MMUART1_DTR_MGPIO12B_OE;
output MMUART1_RI_MGPIO15B_OE;
output MMUART1_RTS_MGPIO11B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI0_SS4_MGPIO19A_OE;
output SPI0_SS5_MGPIO20A_OE;
output SPI0_SS6_MGPIO21A_OE;
output SPI0_SS7_MGPIO22A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module eSRAM_eNVM_access_top_TPSRAM_0_TPSRAM(
       RD_c,
       eSRAM_eNVM_RW_0_ram_wdata,
       eSRAM_eNVM_RW_0_ram_waddr,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       eSRAM_eNVM_RW_0_ram_wen
    );
output [7:0] RD_c;
input  [31:0] eSRAM_eNVM_RW_0_ram_wdata;
input  [4:0] eSRAM_eNVM_RW_0_ram_waddr;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
input  eSRAM_eNVM_RW_0_ram_wen;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    RAM1K18 eSRAM_eNVM_access_top_TPSRAM_0_TPSRAM_R0C0 (.A_DOUT({nc0, 
        nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, nc12, 
        nc13, nc14, nc15, nc16, nc17}), .B_DOUT({nc18, nc19, nc20, 
        nc21, nc22, nc23, nc24, nc25, nc26, nc27, RD_c[7], RD_c[6], 
        RD_c[5], RD_c[4], RD_c[3], RD_c[2], RD_c[1], RD_c[0]}), .BUSY()
        , .A_CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .A_DOUT_CLK(VCC_net_1)
        , .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({
        GND_net_1, VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, 
        eSRAM_eNVM_RW_0_ram_wdata[31], eSRAM_eNVM_RW_0_ram_wdata[30], 
        eSRAM_eNVM_RW_0_ram_wdata[29], eSRAM_eNVM_RW_0_ram_wdata[28], 
        eSRAM_eNVM_RW_0_ram_wdata[27], eSRAM_eNVM_RW_0_ram_wdata[26], 
        eSRAM_eNVM_RW_0_ram_wdata[25], eSRAM_eNVM_RW_0_ram_wdata[24], 
        GND_net_1, eSRAM_eNVM_RW_0_ram_wdata[23], 
        eSRAM_eNVM_RW_0_ram_wdata[22], eSRAM_eNVM_RW_0_ram_wdata[21], 
        eSRAM_eNVM_RW_0_ram_wdata[20], eSRAM_eNVM_RW_0_ram_wdata[19], 
        eSRAM_eNVM_RW_0_ram_wdata[18], eSRAM_eNVM_RW_0_ram_wdata[17], 
        eSRAM_eNVM_RW_0_ram_wdata[16]}), .A_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .A_WEN({VCC_net_1, VCC_net_1}), .B_CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .B_DOUT_CLK(VCC_net_1), 
        .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), .B_BLK({
        eSRAM_eNVM_RW_0_ram_wen, VCC_net_1, VCC_net_1}), 
        .B_DOUT_ARST_N(VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        GND_net_1, eSRAM_eNVM_RW_0_ram_wdata[15], 
        eSRAM_eNVM_RW_0_ram_wdata[14], eSRAM_eNVM_RW_0_ram_wdata[13], 
        eSRAM_eNVM_RW_0_ram_wdata[12], eSRAM_eNVM_RW_0_ram_wdata[11], 
        eSRAM_eNVM_RW_0_ram_wdata[10], eSRAM_eNVM_RW_0_ram_wdata[9], 
        eSRAM_eNVM_RW_0_ram_wdata[8], GND_net_1, 
        eSRAM_eNVM_RW_0_ram_wdata[7], eSRAM_eNVM_RW_0_ram_wdata[6], 
        eSRAM_eNVM_RW_0_ram_wdata[5], eSRAM_eNVM_RW_0_ram_wdata[4], 
        eSRAM_eNVM_RW_0_ram_wdata[3], eSRAM_eNVM_RW_0_ram_wdata[2], 
        eSRAM_eNVM_RW_0_ram_wdata[1], eSRAM_eNVM_RW_0_ram_wdata[0]}), 
        .B_ADDR({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        eSRAM_eNVM_RW_0_ram_waddr[4], eSRAM_eNVM_RW_0_ram_waddr[3], 
        eSRAM_eNVM_RW_0_ram_waddr[2], eSRAM_eNVM_RW_0_ram_waddr[1], 
        eSRAM_eNVM_RW_0_ram_waddr[0], GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .B_WEN({VCC_net_1, VCC_net_1}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, VCC_net_1}), .A_WMODE(GND_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        VCC_net_1}), .B_WMODE(GND_net_1), .SII_LOCK(GND_net_1));
    
endmodule


module eSRAM_eNVM_access_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module CoreResetP_Z6_layer0(
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N,
       FAB_RESET_N_c,
       CORERESETP_0_RESET_N_F2M,
       SYSRESET_POR,
       eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F
    );
output eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
input  eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N;
input  FAB_RESET_N_c;
output CORERESETP_0_RESET_N_F2M;
input  SYSRESET_POR;
input  eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F;

    wire MSS_HPMS_READY_int_net_1, mss_ready_select_net_1, VCC_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        GND_net_1, mss_ready_state_net_1, RESET_N_M2F_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, sm1_areset_n_q1_net_1, 
        sm1_areset_n_clk_base_net_1, POWER_ON_RESET_N_q1_net_1, 
        RESET_N_M2F_q1_net_1, FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        MSS_HPMS_READY_int_4_net_1;
    
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        SYSRESET_POR), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1)
        , .LAT(GND_net_1), .Q(POWER_ON_RESET_N_clk_base_net_1));
    CLKINT MSS_HPMS_READY_int_RNISI68 (.A(MSS_HPMS_READY_int_net_1), 
        .Y(eSRAM_eNVM_access_0_HPMS_READY));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        SYSRESET_POR), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1)
        , .LAT(GND_net_1), .Q(POWER_ON_RESET_N_q1_net_1));
    SLE sm1_areset_n_clk_base (.D(sm1_areset_n_q1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        FAB_RESET_N_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(sm1_areset_n_clk_base_net_1));
    GND GND (.Y(GND_net_1));
    SLE RESET_N_F2M_int (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        sm1_areset_n_clk_base_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(CORERESETP_0_RESET_N_F2M));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_clk_base_net_1));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_q1_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE sm1_areset_n_q1 (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        FAB_RESET_N_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(sm1_areset_n_q1_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(RESET_N_M2F_clk_base_net_1)
        , .ALn(POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(mss_ready_select4_net_1), 
        .ALn(POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_select_net_1));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    
endmodule


module COREAHBLITE_ADDRDEC_Z2_layer0(
       sdec_raw_2,
       AHB_IF_0_BIF_1_HADDR_0,
       AHB_IF_0_BIF_1_HADDR_3,
       masterRegAddrSel
    );
output [0:0] sdec_raw_2;
input  AHB_IF_0_BIF_1_HADDR_0;
input  AHB_IF_0_BIF_1_HADDR_3;
input  masterRegAddrSel;

    wire GND_net_1, VCC_net_1;
    
    CFG3 #( .INIT(8'hCD) )  g0 (.A(AHB_IF_0_BIF_1_HADDR_0), .B(
        masterRegAddrSel), .C(AHB_IF_0_BIF_1_HADDR_3), .Y(
        sdec_raw_2[0]));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module COREAHBLITE_DEFAULTSLAVESM_0s_0_1_0(
       sdec_raw_2,
       AHB_IF_0_BIF_1_HTRANS,
       masterDataInProg,
       SDATASELInt_14,
       SDATASELInt_10,
       SDATASELInt_9,
       SDATASELInt_7,
       SDATASELInt_11,
       SDATASELInt_6,
       SDATASELInt_4,
       SDATASELInt_0,
       SDATASELInt_13,
       SDATASELInt_12,
       SDATASELInt_8,
       SDATASELInt_2,
       defSlaveSMCurrentState,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       defSlaveSMNextState,
       masterRegAddrSel,
       g0_1,
       N_53,
       N_76,
       masterAddrClockEnable,
       N_546,
       CoreAHBLite_0_AHBmslave16_HREADY,
       m0s16DataSel,
       HREADY_M_0_iv_i_0,
       PREVDATASLAVEREADY_iv_i_0
    );
input  [0:0] sdec_raw_2;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
input  [0:0] masterDataInProg;
input  SDATASELInt_14;
input  SDATASELInt_10;
input  SDATASELInt_9;
input  SDATASELInt_7;
input  SDATASELInt_11;
input  SDATASELInt_6;
input  SDATASELInt_4;
input  SDATASELInt_0;
input  SDATASELInt_13;
input  SDATASELInt_12;
input  SDATASELInt_8;
input  SDATASELInt_2;
output defSlaveSMCurrentState;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output defSlaveSMNextState;
input  masterRegAddrSel;
input  g0_1;
output N_53;
input  N_76;
output masterAddrClockEnable;
output N_546;
input  CoreAHBLite_0_AHBmslave16_HREADY;
input  m0s16DataSel;
output HREADY_M_0_iv_i_0;
output PREVDATASLAVEREADY_iv_i_0;

    wire VCC_net_1, GND_net_1, defSlaveSMNextState_0_o2_7_net_1, 
        defSlaveSMNextState_0_o2_8_net_1, 
        defSlaveSMNextState_0_o2_6_net_1, g0_2;
    
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0020) )  defSlaveSMNextState_0_a2_RNIVQFG1 (.A(
        sdec_raw_2[0]), .B(defSlaveSMNextState), .C(
        AHB_IF_0_BIF_1_HTRANS[1]), .D(masterRegAddrSel), .Y(g0_2));
    CFG4 #( .INIT(16'h0F0E) )  defSlaveSMNextState_0_a2 (.A(
        defSlaveSMNextState_0_o2_7_net_1), .B(
        defSlaveSMNextState_0_o2_8_net_1), .C(defSlaveSMCurrentState), 
        .D(defSlaveSMNextState_0_o2_6_net_1), .Y(defSlaveSMNextState));
    SLE defSlaveSMCurrentState_inst_1 (.D(defSlaveSMNextState), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        defSlaveSMCurrentState));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hFFFE) )  defSlaveSMNextState_0_o2_6 (.A(
        SDATASELInt_13), .B(SDATASELInt_12), .C(SDATASELInt_8), .D(
        SDATASELInt_2), .Y(defSlaveSMNextState_0_o2_6_net_1));
    CFG2 #( .INIT(4'h1) )  defSlaveSMNextState_0_a2_RNI6A671 (.A(N_53), 
        .B(defSlaveSMNextState), .Y(HREADY_M_0_iv_i_0));
    CFG4 #( .INIT(16'h1500) )  defSlaveSMNextState_0_o2_RNI2KC11 (.A(
        N_546), .B(CoreAHBLite_0_AHBmslave16_HREADY), .C(
        masterDataInProg[0]), .D(m0s16DataSel), .Y(N_53));
    CFG4 #( .INIT(16'h3200) )  defSlaveSMNextState_0_a2_RNI7NUI5 (.A(
        g0_1), .B(N_53), .C(N_76), .D(g0_2), .Y(masterAddrClockEnable));
    CFG4 #( .INIT(16'hFFFE) )  defSlaveSMNextState_0_o2_7 (.A(
        SDATASELInt_11), .B(SDATASELInt_6), .C(SDATASELInt_4), .D(
        SDATASELInt_0), .Y(defSlaveSMNextState_0_o2_7_net_1));
    CFG3 #( .INIT(8'hFE) )  defSlaveSMNextState_0_o2 (.A(
        defSlaveSMNextState_0_o2_8_net_1), .B(
        defSlaveSMNextState_0_o2_7_net_1), .C(
        defSlaveSMNextState_0_o2_6_net_1), .Y(N_546));
    CFG4 #( .INIT(16'hFFFE) )  defSlaveSMNextState_0_o2_8 (.A(
        SDATASELInt_14), .B(SDATASELInt_10), .C(SDATASELInt_9), .D(
        SDATASELInt_7), .Y(defSlaveSMNextState_0_o2_8_net_1));
    CFG4 #( .INIT(16'h00FB) )  defSlaveSMNextState_0_a2_RNIMUBP (.A(
        N_546), .B(m0s16DataSel), .C(CoreAHBLite_0_AHBmslave16_HREADY), 
        .D(defSlaveSMNextState), .Y(PREVDATASLAVEREADY_iv_i_0));
    
endmodule


module COREAHBLITE_MASTERSTAGE_1_1_85_65536_0s_0_1_0(
       AHB_IF_0_BIF_1_HADDR,
       AHB_IF_0_BIF_1_HTRANS,
       arbRegSMCurrentState_ns_i_0_a2_0_0,
       sdec_raw_2,
       masterDataInProg,
       regHADDR_20,
       regHADDR_21,
       regHADDR_22,
       regHADDR_23,
       regHADDR_24,
       regHADDR_25,
       regHADDR_5,
       regHADDR_6,
       regHADDR_7,
       regHADDR_8,
       regHADDR_9,
       regHADDR_10,
       regHADDR_11,
       regHADDR_12,
       regHADDR_13,
       regHADDR_14,
       regHADDR_15,
       regHADDR_16,
       regHADDR_17,
       regHADDR_18,
       regHADDR_19,
       regHADDR_0,
       regHADDR_1,
       regHADDR_2,
       regHADDR_3,
       regHADDR_4,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       m0s16DataSel,
       m0s16AddrSel_i_0,
       regHWRITE,
       AHB_IF_0_BIF_1_HWRITE,
       regHTRANS,
       masterRegAddrSel,
       N_60,
       N_205,
       N_204,
       N_76,
       defSlaveSMCurrentState,
       defSlaveSMNextState,
       g0_1,
       N_53,
       N_546,
       CoreAHBLite_0_AHBmslave16_HREADY,
       HREADY_M_0_iv_i_0
    );
input  [31:2] AHB_IF_0_BIF_1_HADDR;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
input  [0:0] arbRegSMCurrentState_ns_i_0_a2_0_0;
output [0:0] sdec_raw_2;
input  [0:0] masterDataInProg;
output regHADDR_20;
output regHADDR_21;
output regHADDR_22;
output regHADDR_23;
output regHADDR_24;
output regHADDR_25;
output regHADDR_5;
output regHADDR_6;
output regHADDR_7;
output regHADDR_8;
output regHADDR_9;
output regHADDR_10;
output regHADDR_11;
output regHADDR_12;
output regHADDR_13;
output regHADDR_14;
output regHADDR_15;
output regHADDR_16;
output regHADDR_17;
output regHADDR_18;
output regHADDR_19;
output regHADDR_0;
output regHADDR_1;
output regHADDR_2;
output regHADDR_3;
output regHADDR_4;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output m0s16DataSel;
output m0s16AddrSel_i_0;
output regHWRITE;
input  AHB_IF_0_BIF_1_HWRITE;
output regHTRANS;
output masterRegAddrSel;
input  N_60;
output N_205;
output N_204;
input  N_76;
output defSlaveSMCurrentState;
output defSlaveSMNextState;
input  g0_1;
output N_53;
output N_546;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output HREADY_M_0_iv_i_0;

    wire VCC_net_1, masterAddrClockEnable, GND_net_1, 
        \regHADDR[29]_net_1 , \regHADDR[30]_net_1 , 
        \SDATASELInt[10]_net_1 , \SADDRSEL[10] , 
        PREVDATASLAVEREADY_iv_i_0, \SDATASELInt[11]_net_1 , N_51_i_0, 
        \SDATASELInt[12]_net_1 , \SADDRSEL[12] , 
        \SDATASELInt[13]_net_1 , N_54_i_0, \SDATASELInt[14]_net_1 , 
        \SADDRSEL[14] , \SDATASELInt[15]_net_1 , N_57_i_0, 
        \SDATASELInt[1]_net_1 , \SADDRSEL[1] , \SDATASELInt[3]_net_1 , 
        \SADDRSEL[3] , \SDATASELInt[5]_net_1 , \SADDRSEL[5] , 
        \SDATASELInt[7]_net_1 , \SADDRSEL[7] , \SDATASELInt[8]_net_1 , 
        \SADDRSEL[8] , \SDATASELInt[9]_net_1 , N_48_i_0, 
        d_masterRegAddrSel, N_198, N_264, N_263, N_254;
    
    CFG3 #( .INIT(8'hD8) )  \PREGATEDHADDR_i_m2[29]  (.A(
        masterRegAddrSel), .B(\regHADDR[29]_net_1 ), .C(
        AHB_IF_0_BIF_1_HADDR[29]), .Y(N_205));
    CFG4 #( .INIT(16'hF100) )  masterRegAddrSel_RNIMU0Q1 (.A(
        AHB_IF_0_BIF_1_HADDR[31]), .B(AHB_IF_0_BIF_1_HADDR[28]), .C(
        masterRegAddrSel), .D(N_60), .Y(m0s16AddrSel_i_0));
    SLE \regHADDR[21]  (.D(AHB_IF_0_BIF_1_HADDR[21]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_19));
    SLE \regHADDR[15]  (.D(AHB_IF_0_BIF_1_HADDR[15]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_13));
    SLE \regHADDR[30]  (.D(AHB_IF_0_BIF_1_HADDR[30]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \regHADDR[30]_net_1 ));
    SLE \regHADDR[7]  (.D(AHB_IF_0_BIF_1_HADDR[7]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_5));
    COREAHBLITE_ADDRDEC_Z2_layer0 address_decode (.sdec_raw_2({
        sdec_raw_2[0]}), .AHB_IF_0_BIF_1_HADDR_0(
        AHB_IF_0_BIF_1_HADDR[28]), .AHB_IF_0_BIF_1_HADDR_3(
        AHB_IF_0_BIF_1_HADDR[31]), .masterRegAddrSel(masterRegAddrSel));
    SLE \regHADDR[9]  (.D(AHB_IF_0_BIF_1_HADDR[9]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_7));
    CFG4 #( .INIT(16'h2000) )  \SADDRSEL_0_a2[3]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_263), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[3] ));
    SLE masterRegAddrSel_inst_1 (.D(d_masterRegAddrSel), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        masterRegAddrSel));
    SLE regHTRANS_inst_1 (.D(VCC_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHTRANS));
    CFG3 #( .INIT(8'h01) )  \SDATASELInt_RNO[9]  (.A(N_204), .B(N_205), 
        .C(N_198), .Y(N_48_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0040) )  \SADDRSEL_0_a2[12]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_264), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[12] ));
    SLE \regHADDR[29]  (.D(AHB_IF_0_BIF_1_HADDR[29]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \regHADDR[29]_net_1 ));
    SLE \regHADDR[24]  (.D(AHB_IF_0_BIF_1_HADDR[24]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_22));
    CFG4 #( .INIT(16'h4000) )  \SADDRSEL_0_a2[14]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_264), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[14] ));
    CFG4 #( .INIT(16'h4000) )  \SADDRSEL_0_a2[10]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_263), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[10] ));
    SLE \regHADDR[10]  (.D(AHB_IF_0_BIF_1_HADDR[10]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_8));
    CFG4 #( .INIT(16'h0040) )  \SADDRSEL_0_a2[8]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_263), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[8] ));
    SLE \regHADDR[13]  (.D(AHB_IF_0_BIF_1_HADDR[13]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_11));
    SLE \regHADDR[12]  (.D(AHB_IF_0_BIF_1_HADDR[12]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_10));
    SLE \regHADDR[5]  (.D(AHB_IF_0_BIF_1_HADDR[5]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_3));
    SLE \regHADDR[2]  (.D(AHB_IF_0_BIF_1_HADDR[2]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_0));
    SLE \SDATASELInt[15]  (.D(N_57_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[15]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \SADDRSEL_0_a2_1[8]  (.A(N_204), .B(
        AHB_IF_0_BIF_1_HTRANS[1]), .C(masterRegAddrSel), .Y(N_263));
    SLE \SDATASELInt[14]  (.D(\SADDRSEL[14] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[14]_net_1 ));
    SLE \regHADDR[8]  (.D(AHB_IF_0_BIF_1_HADDR[8]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_6));
    SLE \regHADDR[25]  (.D(AHB_IF_0_BIF_1_HADDR[25]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_23));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h04) )  \SDATASELInt_RNO[11]  (.A(N_204), .B(N_205)
        , .C(N_198), .Y(N_51_i_0));
    SLE \regHADDR[17]  (.D(AHB_IF_0_BIF_1_HADDR[17]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_15));
    CFG3 #( .INIT(8'h08) )  \SADDRSEL_0_a2_1[5]  (.A(N_204), .B(
        AHB_IF_0_BIF_1_HTRANS[1]), .C(masterRegAddrSel), .Y(N_264));
    CFG4 #( .INIT(16'h2000) )  \SADDRSEL_0_a2[7]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_264), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[7] ));
    SLE \regHADDR[6]  (.D(AHB_IF_0_BIF_1_HADDR[6]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_4));
    SLE \regHADDR[16]  (.D(AHB_IF_0_BIF_1_HADDR[16]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_14));
    SLE \SDATASELInt[13]  (.D(N_54_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[13]_net_1 ));
    SLE regHWRITE_inst_1 (.D(AHB_IF_0_BIF_1_HWRITE), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHWRITE));
    SLE \SDATASELInt[9]  (.D(N_48_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[9]_net_1 ));
    SLE \SDATASELInt[1]  (.D(\SADDRSEL[1] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[1]_net_1 ));
    SLE \SDATASELInt[12]  (.D(\SADDRSEL[12] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[12]_net_1 ));
    SLE \regHADDR[11]  (.D(AHB_IF_0_BIF_1_HADDR[11]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_9));
    SLE \SDATASELInt[5]  (.D(\SADDRSEL[5] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[5]_net_1 ));
    CFG2 #( .INIT(4'hE) )  d_masterRegAddrSel_0 (.A(
        masterAddrClockEnable), .B(N_254), .Y(d_masterRegAddrSel));
    SLE \regHADDR[3]  (.D(AHB_IF_0_BIF_1_HADDR[3]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_1));
    CFG4 #( .INIT(16'h0020) )  \SADDRSEL_0_a2[5]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_264), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[5] ));
    SLE \SDATASELInt[3]  (.D(\SADDRSEL[3] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[3]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \SDATASELInt_RNO[15]  (.A(N_204), .B(N_205)
        , .C(N_198), .Y(N_57_i_0));
    SLE \regHADDR[20]  (.D(AHB_IF_0_BIF_1_HADDR[20]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_18));
    SLE \regHADDR[23]  (.D(AHB_IF_0_BIF_1_HADDR[23]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_21));
    SLE \regHADDR[22]  (.D(AHB_IF_0_BIF_1_HADDR[22]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_20));
    CFG3 #( .INIT(8'h02) )  \SDATASELInt_RNO[13]  (.A(N_204), .B(N_205)
        , .C(N_198), .Y(N_54_i_0));
    SLE \SDATASELInt[7]  (.D(\SADDRSEL[7] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[7]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  \SADDRSEL_0_a2[1]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(AHB_IF_0_BIF_1_HADDR[31]), .C(
        N_263), .D(AHB_IF_0_BIF_1_HADDR[29]), .Y(\SADDRSEL[1] ));
    SLE \regHADDR[19]  (.D(AHB_IF_0_BIF_1_HADDR[19]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_17));
    SLE \regHADDR[14]  (.D(AHB_IF_0_BIF_1_HADDR[14]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_12));
    CFG4 #( .INIT(16'hC800) )  d_masterRegAddrSel_0_a2 (.A(N_76), .B(
        masterRegAddrSel), .C(arbRegSMCurrentState_ns_i_0_a2_0_0[0]), 
        .D(m0s16AddrSel_i_0), .Y(N_254));
    CFG4 #( .INIT(16'hDFFF) )  \SADDRSEL_i_o2[9]  (.A(
        AHB_IF_0_BIF_1_HADDR[28]), .B(masterRegAddrSel), .C(
        AHB_IF_0_BIF_1_HTRANS[1]), .D(AHB_IF_0_BIF_1_HADDR[31]), .Y(
        N_198));
    SLE \regHADDR[27]  (.D(AHB_IF_0_BIF_1_HADDR[27]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_25));
    SLE \SDATASELInt[16]  (.D(m0s16AddrSel_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(m0s16DataSel));
    SLE \regHADDR[18]  (.D(AHB_IF_0_BIF_1_HADDR[18]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_16));
    SLE \SDATASELInt[11]  (.D(N_51_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[11]_net_1 ));
    SLE \SDATASELInt[8]  (.D(\SADDRSEL[8] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[8]_net_1 ));
    SLE \regHADDR[4]  (.D(AHB_IF_0_BIF_1_HADDR[4]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_2));
    SLE \regHADDR[26]  (.D(AHB_IF_0_BIF_1_HADDR[26]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(masterAddrClockEnable), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(regHADDR_24));
    SLE \SDATASELInt[10]  (.D(\SADDRSEL[10] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PREVDATASLAVEREADY_iv_i_0), 
        .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDATASELInt[10]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \PREGATEDHADDR_i_m2[30]  (.A(
        masterRegAddrSel), .B(\regHADDR[30]_net_1 ), .C(
        AHB_IF_0_BIF_1_HADDR[30]), .Y(N_204));
    COREAHBLITE_DEFAULTSLAVESM_0s_0_1_0 default_slave_sm (.sdec_raw_2({
        sdec_raw_2[0]}), .AHB_IF_0_BIF_1_HTRANS({
        AHB_IF_0_BIF_1_HTRANS[1]}), .masterDataInProg({
        masterDataInProg[0]}), .SDATASELInt_14(\SDATASELInt[15]_net_1 )
        , .SDATASELInt_10(\SDATASELInt[11]_net_1 ), .SDATASELInt_9(
        \SDATASELInt[10]_net_1 ), .SDATASELInt_7(
        \SDATASELInt[8]_net_1 ), .SDATASELInt_11(
        \SDATASELInt[12]_net_1 ), .SDATASELInt_6(
        \SDATASELInt[7]_net_1 ), .SDATASELInt_4(\SDATASELInt[5]_net_1 )
        , .SDATASELInt_0(\SDATASELInt[1]_net_1 ), .SDATASELInt_13(
        \SDATASELInt[14]_net_1 ), .SDATASELInt_12(
        \SDATASELInt[13]_net_1 ), .SDATASELInt_8(
        \SDATASELInt[9]_net_1 ), .SDATASELInt_2(\SDATASELInt[3]_net_1 )
        , .defSlaveSMCurrentState(defSlaveSMCurrentState), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .defSlaveSMNextState(defSlaveSMNextState), .masterRegAddrSel(
        masterRegAddrSel), .g0_1(g0_1), .N_53(N_53), .N_76(N_76), 
        .masterAddrClockEnable(masterAddrClockEnable), .N_546(N_546), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .m0s16DataSel(m0s16DataSel), 
        .HREADY_M_0_iv_i_0(HREADY_M_0_iv_i_0), 
        .PREVDATASLAVEREADY_iv_i_0(PREVDATASLAVEREADY_iv_i_0));
    
endmodule


module COREAHBLITE_SLAVEARBITER_Z4_layer0_1(
       arbRegSMCurrentState_ns_i_0_a2_0_0,
       sdec_raw_2,
       regHADDR,
       AHB_IF_0_BIF_1_HADDR_26,
       AHB_IF_0_BIF_1_HADDR_29,
       AHB_IF_0_BIF_1_HADDR_25,
       AHB_IF_0_BIF_1_HADDR_24,
       AHB_IF_0_BIF_1_HADDR_23,
       AHB_IF_0_BIF_1_HADDR_22,
       AHB_IF_0_BIF_1_HADDR_21,
       AHB_IF_0_BIF_1_HADDR_20,
       AHB_IF_0_BIF_1_HADDR_19,
       AHB_IF_0_BIF_1_HADDR_18,
       AHB_IF_0_BIF_1_HADDR_17,
       AHB_IF_0_BIF_1_HADDR_16,
       AHB_IF_0_BIF_1_HADDR_15,
       AHB_IF_0_BIF_1_HADDR_14,
       AHB_IF_0_BIF_1_HADDR_13,
       AHB_IF_0_BIF_1_HADDR_12,
       AHB_IF_0_BIF_1_HADDR_11,
       AHB_IF_0_BIF_1_HADDR_10,
       AHB_IF_0_BIF_1_HADDR_9,
       AHB_IF_0_BIF_1_HADDR_8,
       AHB_IF_0_BIF_1_HADDR_7,
       AHB_IF_0_BIF_1_HADDR_6,
       AHB_IF_0_BIF_1_HADDR_5,
       AHB_IF_0_BIF_1_HADDR_4,
       AHB_IF_0_BIF_1_HADDR_3,
       AHB_IF_0_BIF_1_HADDR_2,
       AHB_IF_0_BIF_1_HADDR_1,
       AHB_IF_0_BIF_1_HADDR_0,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       N_60,
       CoreAHBLite_0_AHBmslave16_HREADY,
       N_76,
       m0s16DataSel,
       defSlaveSMNextState,
       N_33_i_0,
       m0s16AddrSel_i_0,
       N_260,
       masterRegAddrSel,
       N_108_i_0,
       regHWRITE,
       AHB_IF_0_BIF_1_HWRITE,
       N_118_i_0,
       regHTRANS,
       N_116_i_0,
       N_114_i_0,
       N_204,
       N_112_i_0,
       N_205,
       N_110_i_0,
       N_39_i_0,
       N_37_i_0,
       N_106_i_0,
       N_104_i_0_0,
       N_102_i_0,
       N_100_i_0,
       N_98_i_0,
       N_96_i_0,
       N_94_i_0,
       N_92_i_0,
       N_90_i_0,
       N_88_i_0,
       N_86_i_0,
       N_17_i_0,
       N_16_i_0,
       N_15_i_0,
       N_78_i_0,
       N_14_i_0,
       N_74_i_0,
       N_72_i_0,
       N_70_i_0,
       N_68_i_0,
       N_13_i_0,
       N_64_i_0,
       N_12_i_0,
       N_11_i_0
    );
output [0:0] arbRegSMCurrentState_ns_i_0_a2_0_0;
input  [0:0] sdec_raw_2;
input  [27:2] regHADDR;
input  AHB_IF_0_BIF_1_HADDR_26;
input  AHB_IF_0_BIF_1_HADDR_29;
input  AHB_IF_0_BIF_1_HADDR_25;
input  AHB_IF_0_BIF_1_HADDR_24;
input  AHB_IF_0_BIF_1_HADDR_23;
input  AHB_IF_0_BIF_1_HADDR_22;
input  AHB_IF_0_BIF_1_HADDR_21;
input  AHB_IF_0_BIF_1_HADDR_20;
input  AHB_IF_0_BIF_1_HADDR_19;
input  AHB_IF_0_BIF_1_HADDR_18;
input  AHB_IF_0_BIF_1_HADDR_17;
input  AHB_IF_0_BIF_1_HADDR_16;
input  AHB_IF_0_BIF_1_HADDR_15;
input  AHB_IF_0_BIF_1_HADDR_14;
input  AHB_IF_0_BIF_1_HADDR_13;
input  AHB_IF_0_BIF_1_HADDR_12;
input  AHB_IF_0_BIF_1_HADDR_11;
input  AHB_IF_0_BIF_1_HADDR_10;
input  AHB_IF_0_BIF_1_HADDR_9;
input  AHB_IF_0_BIF_1_HADDR_8;
input  AHB_IF_0_BIF_1_HADDR_7;
input  AHB_IF_0_BIF_1_HADDR_6;
input  AHB_IF_0_BIF_1_HADDR_5;
input  AHB_IF_0_BIF_1_HADDR_4;
input  AHB_IF_0_BIF_1_HADDR_3;
input  AHB_IF_0_BIF_1_HADDR_2;
input  AHB_IF_0_BIF_1_HADDR_1;
input  AHB_IF_0_BIF_1_HADDR_0;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
input  N_60;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output N_76;
input  m0s16DataSel;
input  defSlaveSMNextState;
output N_33_i_0;
input  m0s16AddrSel_i_0;
output N_260;
input  masterRegAddrSel;
output N_108_i_0;
input  regHWRITE;
input  AHB_IF_0_BIF_1_HWRITE;
output N_118_i_0;
input  regHTRANS;
output N_116_i_0;
output N_114_i_0;
input  N_204;
output N_112_i_0;
input  N_205;
output N_110_i_0;
output N_39_i_0;
output N_37_i_0;
output N_106_i_0;
output N_104_i_0_0;
output N_102_i_0;
output N_100_i_0;
output N_98_i_0;
output N_96_i_0;
output N_94_i_0;
output N_92_i_0;
output N_90_i_0;
output N_88_i_0;
output N_86_i_0;
output N_17_i_0;
output N_16_i_0;
output N_15_i_0;
output N_78_i_0;
output N_14_i_0;
output N_74_i_0;
output N_72_i_0;
output N_70_i_0;
output N_68_i_0;
output N_13_i_0;
output N_64_i_0;
output N_12_i_0;
output N_11_i_0;

    wire \arbRegSMCurrentState[0]_net_1 , VCC_net_1, N_104_i_0, 
        GND_net_1, \arbRegSMCurrentState[1]_net_1 , N_136, 
        \arbRegSMCurrentState[5]_net_1 , N_45_i_0, 
        \arbRegSMCurrentState[9]_net_1 , N_43_i_0, 
        \arbRegSMCurrentState[13]_net_1 , N_41_i_0, N_87, 
        \arbRegSMCurrentState_ns_i_i_a2_1_0[1]_net_1 , N_250;
    
    CFG4 #( .INIT(16'hEEEC) )  \arbRegSMCurrentState_ns_i_i[1]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_250), .C(
        \arbRegSMCurrentState[0]_net_1 ), .D(
        \arbRegSMCurrentState_ns_i_i_a2_1_0[1]_net_1 ), .Y(N_136));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNITNI01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[2]), .D(
        AHB_IF_0_BIF_1_HADDR_0), .Y(N_11_i_0));
    CFG4 #( .INIT(16'hFE00) )  \arbRegSMCurrentState_ns_i_i_a2_1_0[1]  
        (.A(\arbRegSMCurrentState[13]_net_1 ), .B(
        \arbRegSMCurrentState[9]_net_1 ), .C(
        \arbRegSMCurrentState[5]_net_1 ), .D(m0s16AddrSel_i_0), .Y(
        \arbRegSMCurrentState_ns_i_i_a2_1_0[1]_net_1 ));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI987A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[26]), .D(
        AHB_IF_0_BIF_1_HADDR_24), .Y(N_37_i_0));
    CFG4 #( .INIT(16'h0001) )  \arbRegSMCurrentState_RNIFG98[1]  (.A(
        \arbRegSMCurrentState[9]_net_1 ), .B(
        \arbRegSMCurrentState[5]_net_1 ), .C(
        \arbRegSMCurrentState[1]_net_1 ), .D(
        \arbRegSMCurrentState[13]_net_1 ), .Y(N_87));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIVT6A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[21]), .D(
        AHB_IF_0_BIF_1_HADDR_19), .Y(N_98_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI547A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[24]), .D(
        AHB_IF_0_BIF_1_HADDR_22), .Y(N_104_i_0_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI965A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[17]), .D(
        AHB_IF_0_BIF_1_HADDR_15), .Y(N_90_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI327A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[23]), .D(
        AHB_IF_0_BIF_1_HADDR_21), .Y(N_102_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI767A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[25]), .D(
        AHB_IF_0_BIF_1_HADDR_23), .Y(N_106_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI107A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[22]), .D(
        AHB_IF_0_BIF_1_HADDR_20), .Y(N_100_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI9E151[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHWRITE), .D(
        AHB_IF_0_BIF_1_HWRITE), .Y(N_118_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIDA5A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[19]), .D(
        AHB_IF_0_BIF_1_HADDR_17), .Y(N_94_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI1SI01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[4]), .D(
        AHB_IF_0_BIF_1_HADDR_2), .Y(N_64_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNITP4A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[11]), .D(
        AHB_IF_0_BIF_1_HADDR_9), .Y(N_78_i_0));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[0]  (.A(
        CoreAHBLite_0_AHBmslave16_HREADY), .B(N_260), .Y(N_104_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIB6J01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[9]), .D(
        AHB_IF_0_BIF_1_HADDR_7), .Y(N_74_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI3UI01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[5]), .D(
        AHB_IF_0_BIF_1_HADDR_3), .Y(N_13_i_0));
    SLE \arbRegSMCurrentState[0]  (.D(N_104_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[0]_net_1 ));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI745A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[16]), .D(
        AHB_IF_0_BIF_1_HADDR_14), .Y(N_88_i_0));
    CFG3 #( .INIT(8'hB0) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNITQJ11[0]  (.A(regHTRANS), 
        .B(masterRegAddrSel), .C(N_260), .Y(N_116_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI72J01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[7]), .D(
        AHB_IF_0_BIF_1_HADDR_5), .Y(N_70_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIVR4A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[12]), .D(
        AHB_IF_0_BIF_1_HADDR_10), .Y(N_15_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIBA7A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[27]), .D(
        AHB_IF_0_BIF_1_HADDR_25), .Y(N_39_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI50J01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[6]), .D(
        AHB_IF_0_BIF_1_HADDR_4), .Y(N_68_i_0));
    SLE \arbRegSMCurrentState[1]  (.D(N_136), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h8) )  \arbRegSMCurrentState_ns_i_0_a2_RNIH38K[0]  
        (.A(N_260), .B(N_205), .Y(N_110_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNITR6A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[20]), .D(
        AHB_IF_0_BIF_1_HADDR_18), .Y(N_96_i_0));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[13]  (.A(
        m0s16AddrSel_i_0), .B(\arbRegSMCurrentState[13]_net_1 ), .Y(
        N_41_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIRN4A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[10]), .D(
        AHB_IF_0_BIF_1_HADDR_8), .Y(N_14_i_0));
    CFG3 #( .INIT(8'hD0) )  \arbRegSMCurrentState_ns_i_i_a2[1]  (.A(
        m0s16AddrSel_i_0), .B(CoreAHBLite_0_AHBmslave16_HREADY), .C(
        \arbRegSMCurrentState[1]_net_1 ), .Y(N_250));
    CFG2 #( .INIT(4'h8) )  \arbRegSMCurrentState_ns_i_0_a2_RNI9S8K[0]  
        (.A(N_260), .B(N_204), .Y(N_112_i_0));
    CFG3 #( .INIT(8'h31) )  \arbRegSMCurrentState_RNIOAT31[0]  (.A(
        sdec_raw_2[0]), .B(\arbRegSMCurrentState[0]_net_1 ), .C(N_87), 
        .Y(N_76));
    CFG3 #( .INIT(8'h04) )  \arbRegSMCurrentState_RNI988K1[0]  (.A(
        N_76), .B(AHB_IF_0_BIF_1_HADDR_26), .C(masterRegAddrSel), .Y(
        N_108_i_0));
    CFG4 #( .INIT(16'h008C) )  \arbRegSMCurrentState_RNIKBAK2[0]  (.A(
        m0s16DataSel), .B(N_60), .C(defSlaveSMNextState), .D(N_76), .Y(
        N_33_i_0));
    SLE \arbRegSMCurrentState[9]  (.D(N_43_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[9]_net_1 ));
    SLE \arbRegSMCurrentState[13]  (.D(N_41_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[13]_net_1 ));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI525A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[15]), .D(
        AHB_IF_0_BIF_1_HADDR_13), .Y(N_86_i_0));
    CFG3 #( .INIT(8'h37) )  \arbRegSMCurrentState_RNIB5L41[0]  (.A(
        N_60), .B(CoreAHBLite_0_AHBmslave16_HREADY), .C(
        \arbRegSMCurrentState[0]_net_1 ), .Y(
        arbRegSMCurrentState_ns_i_0_a2_0_0[0]));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI94J01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[8]), .D(
        AHB_IF_0_BIF_1_HADDR_6), .Y(N_72_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIB85A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[18]), .D(
        AHB_IF_0_BIF_1_HADDR_16), .Y(N_92_i_0));
    CFG4 #( .INIT(16'hDCCC) )  \arbRegSMCurrentState_ns_i_0_a2[0]  (.A(
        N_87), .B(\arbRegSMCurrentState[0]_net_1 ), .C(sdec_raw_2[0]), 
        .D(N_60), .Y(N_260));
    SLE \arbRegSMCurrentState[5]  (.D(N_45_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \arbRegSMCurrentState[5]_net_1 ));
    CFG3 #( .INIT(8'h08) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNINSVR[0]  (.A(N_260), .B(
        AHB_IF_0_BIF_1_HADDR_29), .C(masterRegAddrSel), .Y(N_114_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNIVPI01[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[3]), .D(
        AHB_IF_0_BIF_1_HADDR_1), .Y(N_12_i_0));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[5]  (.A(
        m0s16AddrSel_i_0), .B(\arbRegSMCurrentState[5]_net_1 ), .Y(
        N_45_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI305A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[14]), .D(
        AHB_IF_0_BIF_1_HADDR_12), .Y(N_17_i_0));
    CFG2 #( .INIT(4'h4) )  \arbRegSMCurrentState_RNO[9]  (.A(
        m0s16AddrSel_i_0), .B(\arbRegSMCurrentState[9]_net_1 ), .Y(
        N_43_i_0));
    CFG4 #( .INIT(16'hC480) )  
        \arbRegSMCurrentState_ns_i_0_a2_RNI1U4A1[0]  (.A(
        masterRegAddrSel), .B(N_260), .C(regHADDR[13]), .D(
        AHB_IF_0_BIF_1_HADDR_11), .Y(N_16_i_0));
    
endmodule


module COREAHBLITE_SLAVESTAGE_0s_0_0_0(
       masterDataInProg,
       AHB_IF_0_BIF_1_HTRANS,
       AHB_IF_0_BIF_1_HWDATA,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       arbRegSMCurrentState_ns_i_0_a2_0_0,
       sdec_raw_2,
       regHADDR,
       AHB_IF_0_BIF_1_HADDR_26,
       AHB_IF_0_BIF_1_HADDR_29,
       AHB_IF_0_BIF_1_HADDR_25,
       AHB_IF_0_BIF_1_HADDR_24,
       AHB_IF_0_BIF_1_HADDR_23,
       AHB_IF_0_BIF_1_HADDR_22,
       AHB_IF_0_BIF_1_HADDR_21,
       AHB_IF_0_BIF_1_HADDR_20,
       AHB_IF_0_BIF_1_HADDR_19,
       AHB_IF_0_BIF_1_HADDR_18,
       AHB_IF_0_BIF_1_HADDR_17,
       AHB_IF_0_BIF_1_HADDR_16,
       AHB_IF_0_BIF_1_HADDR_15,
       AHB_IF_0_BIF_1_HADDR_14,
       AHB_IF_0_BIF_1_HADDR_13,
       AHB_IF_0_BIF_1_HADDR_12,
       AHB_IF_0_BIF_1_HADDR_11,
       AHB_IF_0_BIF_1_HADDR_10,
       AHB_IF_0_BIF_1_HADDR_9,
       AHB_IF_0_BIF_1_HADDR_8,
       AHB_IF_0_BIF_1_HADDR_7,
       AHB_IF_0_BIF_1_HADDR_6,
       AHB_IF_0_BIF_1_HADDR_5,
       AHB_IF_0_BIF_1_HADDR_4,
       AHB_IF_0_BIF_1_HADDR_3,
       AHB_IF_0_BIF_1_HADDR_2,
       AHB_IF_0_BIF_1_HADDR_1,
       AHB_IF_0_BIF_1_HADDR_0,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       N_260,
       CoreAHBLite_0_AHBmslave16_HREADY,
       masterRegAddrSel,
       regHTRANS,
       N_60,
       N_76,
       m0s16DataSel,
       defSlaveSMNextState,
       N_33_i_0,
       m0s16AddrSel_i_0,
       N_108_i_0,
       regHWRITE,
       AHB_IF_0_BIF_1_HWRITE,
       N_118_i_0,
       N_116_i_0,
       N_114_i_0,
       N_204,
       N_112_i_0,
       N_205,
       N_110_i_0,
       N_39_i_0,
       N_37_i_0,
       N_106_i_0,
       N_104_i_0,
       N_102_i_0,
       N_100_i_0,
       N_98_i_0,
       N_96_i_0,
       N_94_i_0,
       N_92_i_0,
       N_90_i_0,
       N_88_i_0,
       N_86_i_0,
       N_17_i_0,
       N_16_i_0,
       N_15_i_0,
       N_78_i_0,
       N_14_i_0,
       N_74_i_0,
       N_72_i_0,
       N_70_i_0,
       N_68_i_0,
       N_13_i_0,
       N_64_i_0,
       N_12_i_0,
       N_11_i_0
    );
output [0:0] masterDataInProg;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
input  [31:0] AHB_IF_0_BIF_1_HWDATA;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
output [0:0] arbRegSMCurrentState_ns_i_0_a2_0_0;
input  [0:0] sdec_raw_2;
input  [27:2] regHADDR;
input  AHB_IF_0_BIF_1_HADDR_26;
input  AHB_IF_0_BIF_1_HADDR_29;
input  AHB_IF_0_BIF_1_HADDR_25;
input  AHB_IF_0_BIF_1_HADDR_24;
input  AHB_IF_0_BIF_1_HADDR_23;
input  AHB_IF_0_BIF_1_HADDR_22;
input  AHB_IF_0_BIF_1_HADDR_21;
input  AHB_IF_0_BIF_1_HADDR_20;
input  AHB_IF_0_BIF_1_HADDR_19;
input  AHB_IF_0_BIF_1_HADDR_18;
input  AHB_IF_0_BIF_1_HADDR_17;
input  AHB_IF_0_BIF_1_HADDR_16;
input  AHB_IF_0_BIF_1_HADDR_15;
input  AHB_IF_0_BIF_1_HADDR_14;
input  AHB_IF_0_BIF_1_HADDR_13;
input  AHB_IF_0_BIF_1_HADDR_12;
input  AHB_IF_0_BIF_1_HADDR_11;
input  AHB_IF_0_BIF_1_HADDR_10;
input  AHB_IF_0_BIF_1_HADDR_9;
input  AHB_IF_0_BIF_1_HADDR_8;
input  AHB_IF_0_BIF_1_HADDR_7;
input  AHB_IF_0_BIF_1_HADDR_6;
input  AHB_IF_0_BIF_1_HADDR_5;
input  AHB_IF_0_BIF_1_HADDR_4;
input  AHB_IF_0_BIF_1_HADDR_3;
input  AHB_IF_0_BIF_1_HADDR_2;
input  AHB_IF_0_BIF_1_HADDR_1;
input  AHB_IF_0_BIF_1_HADDR_0;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output N_260;
input  CoreAHBLite_0_AHBmslave16_HREADY;
input  masterRegAddrSel;
input  regHTRANS;
output N_60;
output N_76;
input  m0s16DataSel;
input  defSlaveSMNextState;
output N_33_i_0;
input  m0s16AddrSel_i_0;
output N_108_i_0;
input  regHWRITE;
input  AHB_IF_0_BIF_1_HWRITE;
output N_118_i_0;
output N_116_i_0;
output N_114_i_0;
input  N_204;
output N_112_i_0;
input  N_205;
output N_110_i_0;
output N_39_i_0;
output N_37_i_0;
output N_106_i_0;
output N_104_i_0;
output N_102_i_0;
output N_100_i_0;
output N_98_i_0;
output N_96_i_0;
output N_94_i_0;
output N_92_i_0;
output N_90_i_0;
output N_88_i_0;
output N_86_i_0;
output N_17_i_0;
output N_16_i_0;
output N_15_i_0;
output N_78_i_0;
output N_14_i_0;
output N_74_i_0;
output N_72_i_0;
output N_70_i_0;
output N_68_i_0;
output N_13_i_0;
output N_64_i_0;
output N_12_i_0;
output N_11_i_0;

    wire VCC_net_1, GND_net_1;
    
    CFG3 #( .INIT(8'hD8) )  g0_1 (.A(masterRegAddrSel), .B(regHTRANS), 
        .C(AHB_IF_0_BIF_1_HTRANS[1]), .Y(N_60));
    CFG2 #( .INIT(4'h8) )  \HWDATA[22]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[22]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[22]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[20]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[20]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[20]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[23]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[23]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[23]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[12]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[12]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[12]));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  \HWDATA[29]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[29]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[29]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[10]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[10]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[10]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[31]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[31]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[31]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[13]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[13]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[13]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[0]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[0]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[0]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[4]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[4]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[4]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[28]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[28]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[28]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[19]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[19]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[19]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[25]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[25]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[25]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[24]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[24]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[24]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[27]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[27]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[27]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[18]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[18]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[18]));
    GND GND (.Y(GND_net_1));
    SLE \masterDataInProg[0]  (.D(N_260), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        CoreAHBLite_0_AHBmslave16_HREADY), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        masterDataInProg[0]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[15]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[15]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[15]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[14]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[14]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[14]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[8]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[8]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[8]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[3]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[3]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[3]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[17]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[17]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[17]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[5]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[5]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[5]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[30]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[30]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[30]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[9]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[9]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[9]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[7]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[7]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[7]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[1]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[1]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[1]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[6]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[6]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[6]));
    COREAHBLITE_SLAVEARBITER_Z4_layer0_1 slave_arbiter (
        .arbRegSMCurrentState_ns_i_0_a2_0_0({
        arbRegSMCurrentState_ns_i_0_a2_0_0[0]}), .sdec_raw_2({
        sdec_raw_2[0]}), .regHADDR({regHADDR[27], regHADDR[26], 
        regHADDR[25], regHADDR[24], regHADDR[23], regHADDR[22], 
        regHADDR[21], regHADDR[20], regHADDR[19], regHADDR[18], 
        regHADDR[17], regHADDR[16], regHADDR[15], regHADDR[14], 
        regHADDR[13], regHADDR[12], regHADDR[11], regHADDR[10], 
        regHADDR[9], regHADDR[8], regHADDR[7], regHADDR[6], 
        regHADDR[5], regHADDR[4], regHADDR[3], regHADDR[2]}), 
        .AHB_IF_0_BIF_1_HADDR_26(AHB_IF_0_BIF_1_HADDR_26), 
        .AHB_IF_0_BIF_1_HADDR_29(AHB_IF_0_BIF_1_HADDR_29), 
        .AHB_IF_0_BIF_1_HADDR_25(AHB_IF_0_BIF_1_HADDR_25), 
        .AHB_IF_0_BIF_1_HADDR_24(AHB_IF_0_BIF_1_HADDR_24), 
        .AHB_IF_0_BIF_1_HADDR_23(AHB_IF_0_BIF_1_HADDR_23), 
        .AHB_IF_0_BIF_1_HADDR_22(AHB_IF_0_BIF_1_HADDR_22), 
        .AHB_IF_0_BIF_1_HADDR_21(AHB_IF_0_BIF_1_HADDR_21), 
        .AHB_IF_0_BIF_1_HADDR_20(AHB_IF_0_BIF_1_HADDR_20), 
        .AHB_IF_0_BIF_1_HADDR_19(AHB_IF_0_BIF_1_HADDR_19), 
        .AHB_IF_0_BIF_1_HADDR_18(AHB_IF_0_BIF_1_HADDR_18), 
        .AHB_IF_0_BIF_1_HADDR_17(AHB_IF_0_BIF_1_HADDR_17), 
        .AHB_IF_0_BIF_1_HADDR_16(AHB_IF_0_BIF_1_HADDR_16), 
        .AHB_IF_0_BIF_1_HADDR_15(AHB_IF_0_BIF_1_HADDR_15), 
        .AHB_IF_0_BIF_1_HADDR_14(AHB_IF_0_BIF_1_HADDR_14), 
        .AHB_IF_0_BIF_1_HADDR_13(AHB_IF_0_BIF_1_HADDR_13), 
        .AHB_IF_0_BIF_1_HADDR_12(AHB_IF_0_BIF_1_HADDR_12), 
        .AHB_IF_0_BIF_1_HADDR_11(AHB_IF_0_BIF_1_HADDR_11), 
        .AHB_IF_0_BIF_1_HADDR_10(AHB_IF_0_BIF_1_HADDR_10), 
        .AHB_IF_0_BIF_1_HADDR_9(AHB_IF_0_BIF_1_HADDR_9), 
        .AHB_IF_0_BIF_1_HADDR_8(AHB_IF_0_BIF_1_HADDR_8), 
        .AHB_IF_0_BIF_1_HADDR_7(AHB_IF_0_BIF_1_HADDR_7), 
        .AHB_IF_0_BIF_1_HADDR_6(AHB_IF_0_BIF_1_HADDR_6), 
        .AHB_IF_0_BIF_1_HADDR_5(AHB_IF_0_BIF_1_HADDR_5), 
        .AHB_IF_0_BIF_1_HADDR_4(AHB_IF_0_BIF_1_HADDR_4), 
        .AHB_IF_0_BIF_1_HADDR_3(AHB_IF_0_BIF_1_HADDR_3), 
        .AHB_IF_0_BIF_1_HADDR_2(AHB_IF_0_BIF_1_HADDR_2), 
        .AHB_IF_0_BIF_1_HADDR_1(AHB_IF_0_BIF_1_HADDR_1), 
        .AHB_IF_0_BIF_1_HADDR_0(AHB_IF_0_BIF_1_HADDR_0), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .N_60(N_60), .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .N_76(N_76), .m0s16DataSel(
        m0s16DataSel), .defSlaveSMNextState(defSlaveSMNextState), 
        .N_33_i_0(N_33_i_0), .m0s16AddrSel_i_0(m0s16AddrSel_i_0), 
        .N_260(N_260), .masterRegAddrSel(masterRegAddrSel), .N_108_i_0(
        N_108_i_0), .regHWRITE(regHWRITE), .AHB_IF_0_BIF_1_HWRITE(
        AHB_IF_0_BIF_1_HWRITE), .N_118_i_0(N_118_i_0), .regHTRANS(
        regHTRANS), .N_116_i_0(N_116_i_0), .N_114_i_0(N_114_i_0), 
        .N_204(N_204), .N_112_i_0(N_112_i_0), .N_205(N_205), 
        .N_110_i_0(N_110_i_0), .N_39_i_0(N_39_i_0), .N_37_i_0(N_37_i_0)
        , .N_106_i_0(N_106_i_0), .N_104_i_0_0(N_104_i_0), .N_102_i_0(
        N_102_i_0), .N_100_i_0(N_100_i_0), .N_98_i_0(N_98_i_0), 
        .N_96_i_0(N_96_i_0), .N_94_i_0(N_94_i_0), .N_92_i_0(N_92_i_0), 
        .N_90_i_0(N_90_i_0), .N_88_i_0(N_88_i_0), .N_86_i_0(N_86_i_0), 
        .N_17_i_0(N_17_i_0), .N_16_i_0(N_16_i_0), .N_15_i_0(N_15_i_0), 
        .N_78_i_0(N_78_i_0), .N_14_i_0(N_14_i_0), .N_74_i_0(N_74_i_0), 
        .N_72_i_0(N_72_i_0), .N_70_i_0(N_70_i_0), .N_68_i_0(N_68_i_0), 
        .N_13_i_0(N_13_i_0), .N_64_i_0(N_64_i_0), .N_12_i_0(N_12_i_0), 
        .N_11_i_0(N_11_i_0));
    CFG2 #( .INIT(4'h8) )  \HWDATA[21]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[21]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[21]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[26]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[26]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[26]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[2]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[2]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[2]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[11]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[11]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[11]));
    CFG2 #( .INIT(4'h8) )  \HWDATA[16]  (.A(masterDataInProg[0]), .B(
        AHB_IF_0_BIF_1_HWDATA[16]), .Y(
        CoreAHBLite_0_AHBmslave16_HWDATA[16]));
    
endmodule


module COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0_0s(
       AHB_IF_0_BIF_1_HADDR,
       AHB_IF_0_BIF_1_HTRANS,
       sdec_raw_2,
       AHB_IF_0_BIF_1_HWDATA,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       m0s16DataSel,
       AHB_IF_0_BIF_1_HWRITE,
       N_60,
       defSlaveSMCurrentState,
       defSlaveSMNextState,
       g0_1,
       N_53,
       N_546,
       CoreAHBLite_0_AHBmslave16_HREADY,
       HREADY_M_0_iv_i_0,
       N_260,
       N_33_i_0,
       N_108_i_0,
       N_118_i_0,
       N_116_i_0,
       N_114_i_0,
       N_112_i_0,
       N_110_i_0,
       N_39_i_0,
       N_37_i_0,
       N_106_i_0,
       N_104_i_0,
       N_102_i_0,
       N_100_i_0,
       N_98_i_0,
       N_96_i_0,
       N_94_i_0,
       N_92_i_0,
       N_90_i_0,
       N_88_i_0,
       N_86_i_0,
       N_17_i_0,
       N_16_i_0,
       N_15_i_0,
       N_78_i_0,
       N_14_i_0,
       N_74_i_0,
       N_72_i_0,
       N_70_i_0,
       N_68_i_0,
       N_13_i_0,
       N_64_i_0,
       N_12_i_0,
       N_11_i_0
    );
input  [31:2] AHB_IF_0_BIF_1_HADDR;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
output [0:0] sdec_raw_2;
input  [31:0] AHB_IF_0_BIF_1_HWDATA;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output m0s16DataSel;
input  AHB_IF_0_BIF_1_HWRITE;
output N_60;
output defSlaveSMCurrentState;
output defSlaveSMNextState;
input  g0_1;
output N_53;
output N_546;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output HREADY_M_0_iv_i_0;
output N_260;
output N_33_i_0;
output N_108_i_0;
output N_118_i_0;
output N_116_i_0;
output N_114_i_0;
output N_112_i_0;
output N_110_i_0;
output N_39_i_0;
output N_37_i_0;
output N_106_i_0;
output N_104_i_0;
output N_102_i_0;
output N_100_i_0;
output N_98_i_0;
output N_96_i_0;
output N_94_i_0;
output N_92_i_0;
output N_90_i_0;
output N_88_i_0;
output N_86_i_0;
output N_17_i_0;
output N_16_i_0;
output N_15_i_0;
output N_78_i_0;
output N_14_i_0;
output N_74_i_0;
output N_72_i_0;
output N_70_i_0;
output N_68_i_0;
output N_13_i_0;
output N_64_i_0;
output N_12_i_0;
output N_11_i_0;

    wire \regHADDR[22] , \regHADDR[23] , \regHADDR[24] , 
        \regHADDR[25] , \regHADDR[26] , \regHADDR[27] , \regHADDR[7] , 
        \regHADDR[8] , \regHADDR[9] , \regHADDR[10] , \regHADDR[11] , 
        \regHADDR[12] , \regHADDR[13] , \regHADDR[14] , \regHADDR[15] , 
        \regHADDR[16] , \regHADDR[17] , \regHADDR[18] , \regHADDR[19] , 
        \regHADDR[20] , \regHADDR[21] , \regHADDR[2] , \regHADDR[3] , 
        \regHADDR[4] , \regHADDR[5] , \regHADDR[6] , 
        \arbRegSMCurrentState_ns_i_0_a2_0_0[0] , \masterDataInProg[0] , 
        m0s16AddrSel_i_0, regHWRITE, regHTRANS, masterRegAddrSel, 
        N_205, N_204, N_76, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    COREAHBLITE_MASTERSTAGE_1_1_85_65536_0s_0_1_0 masterstage_0 (
        .AHB_IF_0_BIF_1_HADDR({AHB_IF_0_BIF_1_HADDR[31], 
        AHB_IF_0_BIF_1_HADDR[30], AHB_IF_0_BIF_1_HADDR[29], 
        AHB_IF_0_BIF_1_HADDR[28], AHB_IF_0_BIF_1_HADDR[27], 
        AHB_IF_0_BIF_1_HADDR[26], AHB_IF_0_BIF_1_HADDR[25], 
        AHB_IF_0_BIF_1_HADDR[24], AHB_IF_0_BIF_1_HADDR[23], 
        AHB_IF_0_BIF_1_HADDR[22], AHB_IF_0_BIF_1_HADDR[21], 
        AHB_IF_0_BIF_1_HADDR[20], AHB_IF_0_BIF_1_HADDR[19], 
        AHB_IF_0_BIF_1_HADDR[18], AHB_IF_0_BIF_1_HADDR[17], 
        AHB_IF_0_BIF_1_HADDR[16], AHB_IF_0_BIF_1_HADDR[15], 
        AHB_IF_0_BIF_1_HADDR[14], AHB_IF_0_BIF_1_HADDR[13], 
        AHB_IF_0_BIF_1_HADDR[12], AHB_IF_0_BIF_1_HADDR[11], 
        AHB_IF_0_BIF_1_HADDR[10], AHB_IF_0_BIF_1_HADDR[9], 
        AHB_IF_0_BIF_1_HADDR[8], AHB_IF_0_BIF_1_HADDR[7], 
        AHB_IF_0_BIF_1_HADDR[6], AHB_IF_0_BIF_1_HADDR[5], 
        AHB_IF_0_BIF_1_HADDR[4], AHB_IF_0_BIF_1_HADDR[3], 
        AHB_IF_0_BIF_1_HADDR[2]}), .AHB_IF_0_BIF_1_HTRANS({
        AHB_IF_0_BIF_1_HTRANS[1]}), 
        .arbRegSMCurrentState_ns_i_0_a2_0_0({
        \arbRegSMCurrentState_ns_i_0_a2_0_0[0] }), .sdec_raw_2({
        sdec_raw_2[0]}), .masterDataInProg({\masterDataInProg[0] }), 
        .regHADDR_20(\regHADDR[22] ), .regHADDR_21(\regHADDR[23] ), 
        .regHADDR_22(\regHADDR[24] ), .regHADDR_23(\regHADDR[25] ), 
        .regHADDR_24(\regHADDR[26] ), .regHADDR_25(\regHADDR[27] ), 
        .regHADDR_5(\regHADDR[7] ), .regHADDR_6(\regHADDR[8] ), 
        .regHADDR_7(\regHADDR[9] ), .regHADDR_8(\regHADDR[10] ), 
        .regHADDR_9(\regHADDR[11] ), .regHADDR_10(\regHADDR[12] ), 
        .regHADDR_11(\regHADDR[13] ), .regHADDR_12(\regHADDR[14] ), 
        .regHADDR_13(\regHADDR[15] ), .regHADDR_14(\regHADDR[16] ), 
        .regHADDR_15(\regHADDR[17] ), .regHADDR_16(\regHADDR[18] ), 
        .regHADDR_17(\regHADDR[19] ), .regHADDR_18(\regHADDR[20] ), 
        .regHADDR_19(\regHADDR[21] ), .regHADDR_0(\regHADDR[2] ), 
        .regHADDR_1(\regHADDR[3] ), .regHADDR_2(\regHADDR[4] ), 
        .regHADDR_3(\regHADDR[5] ), .regHADDR_4(\regHADDR[6] ), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .m0s16DataSel(m0s16DataSel), .m0s16AddrSel_i_0(
        m0s16AddrSel_i_0), .regHWRITE(regHWRITE), 
        .AHB_IF_0_BIF_1_HWRITE(AHB_IF_0_BIF_1_HWRITE), .regHTRANS(
        regHTRANS), .masterRegAddrSel(masterRegAddrSel), .N_60(N_60), 
        .N_205(N_205), .N_204(N_204), .N_76(N_76), 
        .defSlaveSMCurrentState(defSlaveSMCurrentState), 
        .defSlaveSMNextState(defSlaveSMNextState), .g0_1(g0_1), .N_53(
        N_53), .N_546(N_546), .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .HREADY_M_0_iv_i_0(
        HREADY_M_0_iv_i_0));
    COREAHBLITE_SLAVESTAGE_0s_0_0_0 slavestage_16 (.masterDataInProg({
        \masterDataInProg[0] }), .AHB_IF_0_BIF_1_HTRANS({
        AHB_IF_0_BIF_1_HTRANS[1]}), .AHB_IF_0_BIF_1_HWDATA({
        AHB_IF_0_BIF_1_HWDATA[31], AHB_IF_0_BIF_1_HWDATA[30], 
        AHB_IF_0_BIF_1_HWDATA[29], AHB_IF_0_BIF_1_HWDATA[28], 
        AHB_IF_0_BIF_1_HWDATA[27], AHB_IF_0_BIF_1_HWDATA[26], 
        AHB_IF_0_BIF_1_HWDATA[25], AHB_IF_0_BIF_1_HWDATA[24], 
        AHB_IF_0_BIF_1_HWDATA[23], AHB_IF_0_BIF_1_HWDATA[22], 
        AHB_IF_0_BIF_1_HWDATA[21], AHB_IF_0_BIF_1_HWDATA[20], 
        AHB_IF_0_BIF_1_HWDATA[19], AHB_IF_0_BIF_1_HWDATA[18], 
        AHB_IF_0_BIF_1_HWDATA[17], AHB_IF_0_BIF_1_HWDATA[16], 
        AHB_IF_0_BIF_1_HWDATA[15], AHB_IF_0_BIF_1_HWDATA[14], 
        AHB_IF_0_BIF_1_HWDATA[13], AHB_IF_0_BIF_1_HWDATA[12], 
        AHB_IF_0_BIF_1_HWDATA[11], AHB_IF_0_BIF_1_HWDATA[10], 
        AHB_IF_0_BIF_1_HWDATA[9], AHB_IF_0_BIF_1_HWDATA[8], 
        AHB_IF_0_BIF_1_HWDATA[7], AHB_IF_0_BIF_1_HWDATA[6], 
        AHB_IF_0_BIF_1_HWDATA[5], AHB_IF_0_BIF_1_HWDATA[4], 
        AHB_IF_0_BIF_1_HWDATA[3], AHB_IF_0_BIF_1_HWDATA[2], 
        AHB_IF_0_BIF_1_HWDATA[1], AHB_IF_0_BIF_1_HWDATA[0]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), 
        .arbRegSMCurrentState_ns_i_0_a2_0_0({
        \arbRegSMCurrentState_ns_i_0_a2_0_0[0] }), .sdec_raw_2({
        sdec_raw_2[0]}), .regHADDR({\regHADDR[27] , \regHADDR[26] , 
        \regHADDR[25] , \regHADDR[24] , \regHADDR[23] , \regHADDR[22] , 
        \regHADDR[21] , \regHADDR[20] , \regHADDR[19] , \regHADDR[18] , 
        \regHADDR[17] , \regHADDR[16] , \regHADDR[15] , \regHADDR[14] , 
        \regHADDR[13] , \regHADDR[12] , \regHADDR[11] , \regHADDR[10] , 
        \regHADDR[9] , \regHADDR[8] , \regHADDR[7] , \regHADDR[6] , 
        \regHADDR[5] , \regHADDR[4] , \regHADDR[3] , \regHADDR[2] }), 
        .AHB_IF_0_BIF_1_HADDR_26(AHB_IF_0_BIF_1_HADDR[28]), 
        .AHB_IF_0_BIF_1_HADDR_29(AHB_IF_0_BIF_1_HADDR[31]), 
        .AHB_IF_0_BIF_1_HADDR_25(AHB_IF_0_BIF_1_HADDR[27]), 
        .AHB_IF_0_BIF_1_HADDR_24(AHB_IF_0_BIF_1_HADDR[26]), 
        .AHB_IF_0_BIF_1_HADDR_23(AHB_IF_0_BIF_1_HADDR[25]), 
        .AHB_IF_0_BIF_1_HADDR_22(AHB_IF_0_BIF_1_HADDR[24]), 
        .AHB_IF_0_BIF_1_HADDR_21(AHB_IF_0_BIF_1_HADDR[23]), 
        .AHB_IF_0_BIF_1_HADDR_20(AHB_IF_0_BIF_1_HADDR[22]), 
        .AHB_IF_0_BIF_1_HADDR_19(AHB_IF_0_BIF_1_HADDR[21]), 
        .AHB_IF_0_BIF_1_HADDR_18(AHB_IF_0_BIF_1_HADDR[20]), 
        .AHB_IF_0_BIF_1_HADDR_17(AHB_IF_0_BIF_1_HADDR[19]), 
        .AHB_IF_0_BIF_1_HADDR_16(AHB_IF_0_BIF_1_HADDR[18]), 
        .AHB_IF_0_BIF_1_HADDR_15(AHB_IF_0_BIF_1_HADDR[17]), 
        .AHB_IF_0_BIF_1_HADDR_14(AHB_IF_0_BIF_1_HADDR[16]), 
        .AHB_IF_0_BIF_1_HADDR_13(AHB_IF_0_BIF_1_HADDR[15]), 
        .AHB_IF_0_BIF_1_HADDR_12(AHB_IF_0_BIF_1_HADDR[14]), 
        .AHB_IF_0_BIF_1_HADDR_11(AHB_IF_0_BIF_1_HADDR[13]), 
        .AHB_IF_0_BIF_1_HADDR_10(AHB_IF_0_BIF_1_HADDR[12]), 
        .AHB_IF_0_BIF_1_HADDR_9(AHB_IF_0_BIF_1_HADDR[11]), 
        .AHB_IF_0_BIF_1_HADDR_8(AHB_IF_0_BIF_1_HADDR[10]), 
        .AHB_IF_0_BIF_1_HADDR_7(AHB_IF_0_BIF_1_HADDR[9]), 
        .AHB_IF_0_BIF_1_HADDR_6(AHB_IF_0_BIF_1_HADDR[8]), 
        .AHB_IF_0_BIF_1_HADDR_5(AHB_IF_0_BIF_1_HADDR[7]), 
        .AHB_IF_0_BIF_1_HADDR_4(AHB_IF_0_BIF_1_HADDR[6]), 
        .AHB_IF_0_BIF_1_HADDR_3(AHB_IF_0_BIF_1_HADDR[5]), 
        .AHB_IF_0_BIF_1_HADDR_2(AHB_IF_0_BIF_1_HADDR[4]), 
        .AHB_IF_0_BIF_1_HADDR_1(AHB_IF_0_BIF_1_HADDR[3]), 
        .AHB_IF_0_BIF_1_HADDR_0(AHB_IF_0_BIF_1_HADDR[2]), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .N_260(N_260), .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .masterRegAddrSel(
        masterRegAddrSel), .regHTRANS(regHTRANS), .N_60(N_60), .N_76(
        N_76), .m0s16DataSel(m0s16DataSel), .defSlaveSMNextState(
        defSlaveSMNextState), .N_33_i_0(N_33_i_0), .m0s16AddrSel_i_0(
        m0s16AddrSel_i_0), .N_108_i_0(N_108_i_0), .regHWRITE(regHWRITE)
        , .AHB_IF_0_BIF_1_HWRITE(AHB_IF_0_BIF_1_HWRITE), .N_118_i_0(
        N_118_i_0), .N_116_i_0(N_116_i_0), .N_114_i_0(N_114_i_0), 
        .N_204(N_204), .N_112_i_0(N_112_i_0), .N_205(N_205), 
        .N_110_i_0(N_110_i_0), .N_39_i_0(N_39_i_0), .N_37_i_0(N_37_i_0)
        , .N_106_i_0(N_106_i_0), .N_104_i_0(N_104_i_0), .N_102_i_0(
        N_102_i_0), .N_100_i_0(N_100_i_0), .N_98_i_0(N_98_i_0), 
        .N_96_i_0(N_96_i_0), .N_94_i_0(N_94_i_0), .N_92_i_0(N_92_i_0), 
        .N_90_i_0(N_90_i_0), .N_88_i_0(N_88_i_0), .N_86_i_0(N_86_i_0), 
        .N_17_i_0(N_17_i_0), .N_16_i_0(N_16_i_0), .N_15_i_0(N_15_i_0), 
        .N_78_i_0(N_78_i_0), .N_14_i_0(N_14_i_0), .N_74_i_0(N_74_i_0), 
        .N_72_i_0(N_72_i_0), .N_70_i_0(N_70_i_0), .N_68_i_0(N_68_i_0), 
        .N_13_i_0(N_13_i_0), .N_64_i_0(N_64_i_0), .N_12_i_0(N_12_i_0), 
        .N_11_i_0(N_11_i_0));
    
endmodule


module CoreAHBLite_Z5_layer0(
       AHB_IF_0_BIF_1_HADDR,
       AHB_IF_0_BIF_1_HTRANS,
       sdec_raw_2,
       AHB_IF_0_BIF_1_HWDATA,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       m0s16DataSel,
       AHB_IF_0_BIF_1_HWRITE,
       N_60,
       defSlaveSMCurrentState,
       defSlaveSMNextState,
       g0_1,
       N_53,
       N_546,
       CoreAHBLite_0_AHBmslave16_HREADY,
       HREADY_M_0_iv_i_0,
       N_260,
       N_33_i_0,
       N_108_i_0,
       N_118_i_0,
       N_116_i_0,
       N_114_i_0,
       N_112_i_0,
       N_110_i_0,
       N_39_i_0,
       N_37_i_0,
       N_106_i_0,
       N_104_i_0,
       N_102_i_0,
       N_100_i_0,
       N_98_i_0,
       N_96_i_0,
       N_94_i_0,
       N_92_i_0,
       N_90_i_0,
       N_88_i_0,
       N_86_i_0,
       N_17_i_0,
       N_16_i_0,
       N_15_i_0,
       N_78_i_0,
       N_14_i_0,
       N_74_i_0,
       N_72_i_0,
       N_70_i_0,
       N_68_i_0,
       N_13_i_0,
       N_64_i_0,
       N_12_i_0,
       N_11_i_0
    );
input  [31:2] AHB_IF_0_BIF_1_HADDR;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
output [0:0] sdec_raw_2;
input  [31:0] AHB_IF_0_BIF_1_HWDATA;
output [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output m0s16DataSel;
input  AHB_IF_0_BIF_1_HWRITE;
output N_60;
output defSlaveSMCurrentState;
output defSlaveSMNextState;
input  g0_1;
output N_53;
output N_546;
input  CoreAHBLite_0_AHBmslave16_HREADY;
output HREADY_M_0_iv_i_0;
output N_260;
output N_33_i_0;
output N_108_i_0;
output N_118_i_0;
output N_116_i_0;
output N_114_i_0;
output N_112_i_0;
output N_110_i_0;
output N_39_i_0;
output N_37_i_0;
output N_106_i_0;
output N_104_i_0;
output N_102_i_0;
output N_100_i_0;
output N_98_i_0;
output N_96_i_0;
output N_94_i_0;
output N_92_i_0;
output N_90_i_0;
output N_88_i_0;
output N_86_i_0;
output N_17_i_0;
output N_16_i_0;
output N_15_i_0;
output N_78_i_0;
output N_14_i_0;
output N_74_i_0;
output N_72_i_0;
output N_70_i_0;
output N_68_i_0;
output N_13_i_0;
output N_64_i_0;
output N_12_i_0;
output N_11_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    COREAHBLITE_MATRIX4X16_1_1_85_65536_0_0_0_0s matrix4x16 (
        .AHB_IF_0_BIF_1_HADDR({AHB_IF_0_BIF_1_HADDR[31], 
        AHB_IF_0_BIF_1_HADDR[30], AHB_IF_0_BIF_1_HADDR[29], 
        AHB_IF_0_BIF_1_HADDR[28], AHB_IF_0_BIF_1_HADDR[27], 
        AHB_IF_0_BIF_1_HADDR[26], AHB_IF_0_BIF_1_HADDR[25], 
        AHB_IF_0_BIF_1_HADDR[24], AHB_IF_0_BIF_1_HADDR[23], 
        AHB_IF_0_BIF_1_HADDR[22], AHB_IF_0_BIF_1_HADDR[21], 
        AHB_IF_0_BIF_1_HADDR[20], AHB_IF_0_BIF_1_HADDR[19], 
        AHB_IF_0_BIF_1_HADDR[18], AHB_IF_0_BIF_1_HADDR[17], 
        AHB_IF_0_BIF_1_HADDR[16], AHB_IF_0_BIF_1_HADDR[15], 
        AHB_IF_0_BIF_1_HADDR[14], AHB_IF_0_BIF_1_HADDR[13], 
        AHB_IF_0_BIF_1_HADDR[12], AHB_IF_0_BIF_1_HADDR[11], 
        AHB_IF_0_BIF_1_HADDR[10], AHB_IF_0_BIF_1_HADDR[9], 
        AHB_IF_0_BIF_1_HADDR[8], AHB_IF_0_BIF_1_HADDR[7], 
        AHB_IF_0_BIF_1_HADDR[6], AHB_IF_0_BIF_1_HADDR[5], 
        AHB_IF_0_BIF_1_HADDR[4], AHB_IF_0_BIF_1_HADDR[3], 
        AHB_IF_0_BIF_1_HADDR[2]}), .AHB_IF_0_BIF_1_HTRANS({
        AHB_IF_0_BIF_1_HTRANS[1]}), .sdec_raw_2({sdec_raw_2[0]}), 
        .AHB_IF_0_BIF_1_HWDATA({AHB_IF_0_BIF_1_HWDATA[31], 
        AHB_IF_0_BIF_1_HWDATA[30], AHB_IF_0_BIF_1_HWDATA[29], 
        AHB_IF_0_BIF_1_HWDATA[28], AHB_IF_0_BIF_1_HWDATA[27], 
        AHB_IF_0_BIF_1_HWDATA[26], AHB_IF_0_BIF_1_HWDATA[25], 
        AHB_IF_0_BIF_1_HWDATA[24], AHB_IF_0_BIF_1_HWDATA[23], 
        AHB_IF_0_BIF_1_HWDATA[22], AHB_IF_0_BIF_1_HWDATA[21], 
        AHB_IF_0_BIF_1_HWDATA[20], AHB_IF_0_BIF_1_HWDATA[19], 
        AHB_IF_0_BIF_1_HWDATA[18], AHB_IF_0_BIF_1_HWDATA[17], 
        AHB_IF_0_BIF_1_HWDATA[16], AHB_IF_0_BIF_1_HWDATA[15], 
        AHB_IF_0_BIF_1_HWDATA[14], AHB_IF_0_BIF_1_HWDATA[13], 
        AHB_IF_0_BIF_1_HWDATA[12], AHB_IF_0_BIF_1_HWDATA[11], 
        AHB_IF_0_BIF_1_HWDATA[10], AHB_IF_0_BIF_1_HWDATA[9], 
        AHB_IF_0_BIF_1_HWDATA[8], AHB_IF_0_BIF_1_HWDATA[7], 
        AHB_IF_0_BIF_1_HWDATA[6], AHB_IF_0_BIF_1_HWDATA[5], 
        AHB_IF_0_BIF_1_HWDATA[4], AHB_IF_0_BIF_1_HWDATA[3], 
        AHB_IF_0_BIF_1_HWDATA[2], AHB_IF_0_BIF_1_HWDATA[1], 
        AHB_IF_0_BIF_1_HWDATA[0]}), .CoreAHBLite_0_AHBmslave16_HWDATA({
        CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .m0s16DataSel(m0s16DataSel), .AHB_IF_0_BIF_1_HWRITE(
        AHB_IF_0_BIF_1_HWRITE), .N_60(N_60), .defSlaveSMCurrentState(
        defSlaveSMCurrentState), .defSlaveSMNextState(
        defSlaveSMNextState), .g0_1(g0_1), .N_53(N_53), .N_546(N_546), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .HREADY_M_0_iv_i_0(
        HREADY_M_0_iv_i_0), .N_260(N_260), .N_33_i_0(N_33_i_0), 
        .N_108_i_0(N_108_i_0), .N_118_i_0(N_118_i_0), .N_116_i_0(
        N_116_i_0), .N_114_i_0(N_114_i_0), .N_112_i_0(N_112_i_0), 
        .N_110_i_0(N_110_i_0), .N_39_i_0(N_39_i_0), .N_37_i_0(N_37_i_0)
        , .N_106_i_0(N_106_i_0), .N_104_i_0(N_104_i_0), .N_102_i_0(
        N_102_i_0), .N_100_i_0(N_100_i_0), .N_98_i_0(N_98_i_0), 
        .N_96_i_0(N_96_i_0), .N_94_i_0(N_94_i_0), .N_92_i_0(N_92_i_0), 
        .N_90_i_0(N_90_i_0), .N_88_i_0(N_88_i_0), .N_86_i_0(N_86_i_0), 
        .N_17_i_0(N_17_i_0), .N_16_i_0(N_16_i_0), .N_15_i_0(N_15_i_0), 
        .N_78_i_0(N_78_i_0), .N_14_i_0(N_14_i_0), .N_74_i_0(N_74_i_0), 
        .N_72_i_0(N_72_i_0), .N_70_i_0(N_70_i_0), .N_68_i_0(N_68_i_0), 
        .N_13_i_0(N_13_i_0), .N_64_i_0(N_64_i_0), .N_12_i_0(N_12_i_0), 
        .N_11_i_0(N_11_i_0));
    GND GND (.Y(GND_net_1));
    
endmodule


module eSRAM_eNVM_access_CCC_0_FCCC(
       eSRAM_eNVM_access_0_FIC_0_CLK,
       LOCK,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output eSRAM_eNVM_access_0_FIC_0_CLK;
output LOCK;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST (.A(GL0_net), .Y(eSRAM_eNVM_access_0_FIC_0_CLK));
    CCC #( .INIT(210'h0000007FB8000044D64000318C6318C1F18C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(LOCK), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module eSRAM_eNVM_access_HPMS(
       sdec_raw_2,
       AHB_IF_0_BIF_1_HRDATA,
       CoreAHBLite_0_AHBmslave16_HWDATA,
       N_60,
       CoreAHBLite_0_AHBmslave16_HREADY,
       g0_1,
       N_546,
       m0s16DataSel,
       eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N,
       eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F,
       N_11_i_0,
       N_12_i_0,
       N_64_i_0,
       N_13_i_0,
       N_68_i_0,
       N_70_i_0,
       N_72_i_0,
       N_74_i_0,
       N_14_i_0,
       N_78_i_0,
       N_15_i_0,
       N_16_i_0,
       N_17_i_0,
       N_86_i_0,
       N_88_i_0,
       N_90_i_0,
       N_92_i_0,
       N_94_i_0,
       N_96_i_0,
       N_98_i_0,
       N_100_i_0,
       N_102_i_0,
       N_104_i_0,
       N_106_i_0,
       N_37_i_0,
       N_39_i_0,
       N_108_i_0,
       N_110_i_0,
       N_112_i_0,
       N_114_i_0,
       N_260,
       N_116_i_0,
       N_33_i_0,
       N_118_i_0,
       LOCK,
       CORERESETP_0_RESET_N_F2M,
       eSRAM_eNVM_access_0_FIC_0_CLK
    );
input  [0:0] sdec_raw_2;
output [31:0] AHB_IF_0_BIF_1_HRDATA;
input  [31:0] CoreAHBLite_0_AHBmslave16_HWDATA;
input  N_60;
inout  CoreAHBLite_0_AHBmslave16_HREADY;
output g0_1;
input  N_546;
input  m0s16DataSel;
output eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N;
output eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F;
input  N_11_i_0;
input  N_12_i_0;
input  N_64_i_0;
input  N_13_i_0;
input  N_68_i_0;
input  N_70_i_0;
input  N_72_i_0;
input  N_74_i_0;
input  N_14_i_0;
input  N_78_i_0;
input  N_15_i_0;
input  N_16_i_0;
input  N_17_i_0;
input  N_86_i_0;
input  N_88_i_0;
input  N_90_i_0;
input  N_92_i_0;
input  N_94_i_0;
input  N_96_i_0;
input  N_98_i_0;
input  N_100_i_0;
input  N_102_i_0;
input  N_104_i_0;
input  N_106_i_0;
input  N_37_i_0;
input  N_39_i_0;
input  N_108_i_0;
input  N_110_i_0;
input  N_112_i_0;
input  N_114_i_0;
input  N_260;
input  N_116_i_0;
input  N_33_i_0;
input  N_118_i_0;
input  LOCK;
input  CORERESETP_0_RESET_N_F2M;
input  eSRAM_eNVM_access_0_FIC_0_CLK;

    wire \CoreAHBLite_0_AHBmslave16_HRDATA[0] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[31] , VCC_net_1, GND_net_1;
    
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_4 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[5] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[5]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_16 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[17] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[17]));
    CFG3 #( .INIT(8'h7F) )  MSS_ADLIB_INST_RNIET4T1 (.A(N_60), .B(
        sdec_raw_2[0]), .C(CoreAHBLite_0_AHBmslave16_HREADY), .Y(g0_1));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_3 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[4] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[4]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_27 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[28] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[28]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_14 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[15] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[15]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_11 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[12] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[12]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_0 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[1] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[1]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_26 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[27] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[27]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_9 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[10] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[10]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_19 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[20] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[20]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_18 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[19] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[19]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_13 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[14] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[14]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_24 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[25] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[25]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_12 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[13] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[13]));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[0] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[0]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_10 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[11] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[11]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_15 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[16] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[16]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_21 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[22] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[22]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_29 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[30] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[30]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_28 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[29] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[29]));
    MSS_025 #( .INIT(1438'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE400000000000010000000000F11C000001FEDFFC010842108421000001FE34001FF8000000000000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(100.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({\CoreAHBLite_0_AHBmslave16_HRDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HRDATA[0] }), .F_FM0_READYOUT(
        CoreAHBLite_0_AHBmslave16_HREADY), .F_FM0_RESP(), .F_HM0_ADDR({
        nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, 
        nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, 
        nc29, nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, 
        nc39}), .F_HM0_ENABLE(), .F_HM0_SEL(), .F_HM0_SIZE({nc40, nc41})
        , .F_HM0_TRANS1(), .F_HM0_WDATA({nc42, nc43, nc44, nc45, nc46, 
        nc47, nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, nc56, 
        nc57, nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, 
        nc67, nc68, nc69, nc70, nc71, nc72, nc73}), .F_HM0_WRITE(), 
        .FAB_CHRGVBUS(), .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), 
        .FAB_DPPULLDOWN(), .FAB_DRVVBUS(), .FAB_IDPULLUP(), 
        .FAB_OPMODE({nc74, nc75}), .FAB_SUSPENDM(), .FAB_TERMSEL(), 
        .FAB_TXVALID(), .FAB_VCONTROL({nc76, nc77, nc78, nc79}), 
        .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({nc80, nc81}), 
        .FAB_XDATAOUT({nc82, nc83, nc84, nc85, nc86, nc87, nc88, nc89})
        , .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc90, nc91}), 
        .FIC32_1_MASTER({nc92, nc93}), .FPGA_RESET_N(
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), 
        .H2F_INTERRUPT({nc94, nc95, nc96, nc97, nc98, nc99, nc100, 
        nc101, nc102, nc103, nc104, nc105, nc106, nc107, nc108, nc109})
        , .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc110, nc111, nc112, nc113, nc114, nc115, 
        nc116, nc117, nc118, nc119, nc120, nc121, nc122, nc123}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc124, nc125, nc126, nc127, nc128, nc129, 
        nc130, nc131, nc132, nc133, nc134, nc135, nc136, nc137, nc138, 
        nc139, nc140, nc141, nc142, nc143, nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, nc151, nc152, nc153, nc154, nc155}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc156, nc157, nc158, nc159, 
        nc160, nc161, nc162, nc163, nc164, nc165}), .TRACECLK(), 
        .TRACEDATA({nc166, nc167, nc168, nc169}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc170, nc171, nc172, 
        nc173}), .TXDF({nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc182, nc183, nc184, nc185})
        , .F_BRESP_HRESP0({nc186, nc187}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc188, nc189, nc190, nc191, nc192, nc193, 
        nc194, nc195, nc196, nc197, nc198, nc199, nc200, nc201, nc202, 
        nc203, nc204, nc205, nc206, nc207, nc208, nc209, nc210, nc211, 
        nc212, nc213, nc214, nc215, nc216, nc217, nc218, nc219, nc220, 
        nc221, nc222, nc223, nc224, nc225, nc226, nc227, nc228, nc229, 
        nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, nc238, 
        nc239, nc240, nc241, nc242, nc243, nc244, nc245, nc246, nc247, 
        nc248, nc249, nc250, nc251}), .F_RID({nc252, nc253, nc254, 
        nc255}), .F_RLAST(), .F_RRESP_HRESP1({nc256, nc257}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc258, nc259, 
        nc260, nc261, nc262, nc263, nc264, nc265, nc266, nc267, nc268, 
        nc269, nc270, nc271, nc272, nc273}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(VCC_net_1), 
        .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({N_114_i_0, 
        N_112_i_0, N_110_i_0, N_108_i_0, N_39_i_0, N_37_i_0, N_106_i_0, 
        N_104_i_0, N_102_i_0, N_100_i_0, N_98_i_0, N_96_i_0, N_94_i_0, 
        N_92_i_0, N_90_i_0, N_88_i_0, N_86_i_0, N_17_i_0, N_16_i_0, 
        N_15_i_0, N_78_i_0, N_14_i_0, N_74_i_0, N_72_i_0, N_70_i_0, 
        N_68_i_0, N_13_i_0, N_64_i_0, N_12_i_0, N_11_i_0, GND_net_1, 
        GND_net_1}), .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(
        GND_net_1), .F_FM0_READY(CoreAHBLite_0_AHBmslave16_HREADY), 
        .F_FM0_SEL(N_260), .F_FM0_SIZE({N_116_i_0, GND_net_1}), 
        .F_FM0_TRANS1(N_33_i_0), .F_FM0_WDATA({
        CoreAHBLite_0_AHBmslave16_HWDATA[31], 
        CoreAHBLite_0_AHBmslave16_HWDATA[30], 
        CoreAHBLite_0_AHBmslave16_HWDATA[29], 
        CoreAHBLite_0_AHBmslave16_HWDATA[28], 
        CoreAHBLite_0_AHBmslave16_HWDATA[27], 
        CoreAHBLite_0_AHBmslave16_HWDATA[26], 
        CoreAHBLite_0_AHBmslave16_HWDATA[25], 
        CoreAHBLite_0_AHBmslave16_HWDATA[24], 
        CoreAHBLite_0_AHBmslave16_HWDATA[23], 
        CoreAHBLite_0_AHBmslave16_HWDATA[22], 
        CoreAHBLite_0_AHBmslave16_HWDATA[21], 
        CoreAHBLite_0_AHBmslave16_HWDATA[20], 
        CoreAHBLite_0_AHBmslave16_HWDATA[19], 
        CoreAHBLite_0_AHBmslave16_HWDATA[18], 
        CoreAHBLite_0_AHBmslave16_HWDATA[17], 
        CoreAHBLite_0_AHBmslave16_HWDATA[16], 
        CoreAHBLite_0_AHBmslave16_HWDATA[15], 
        CoreAHBLite_0_AHBmslave16_HWDATA[14], 
        CoreAHBLite_0_AHBmslave16_HWDATA[13], 
        CoreAHBLite_0_AHBmslave16_HWDATA[12], 
        CoreAHBLite_0_AHBmslave16_HWDATA[11], 
        CoreAHBLite_0_AHBmslave16_HWDATA[10], 
        CoreAHBLite_0_AHBmslave16_HWDATA[9], 
        CoreAHBLite_0_AHBmslave16_HWDATA[8], 
        CoreAHBLite_0_AHBmslave16_HWDATA[7], 
        CoreAHBLite_0_AHBmslave16_HWDATA[6], 
        CoreAHBLite_0_AHBmslave16_HWDATA[5], 
        CoreAHBLite_0_AHBmslave16_HWDATA[4], 
        CoreAHBLite_0_AHBmslave16_HWDATA[3], 
        CoreAHBLite_0_AHBmslave16_HWDATA[2], 
        CoreAHBLite_0_AHBmslave16_HWDATA[1], 
        CoreAHBLite_0_AHBmslave16_HWDATA[0]}), .F_FM0_WRITE(N_118_i_0), 
        .F_HM0_RDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F_HM0_READY(VCC_net_1), 
        .F_HM0_RESP(GND_net_1), .FAB_AVALID(VCC_net_1), 
        .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        GND_net_1), .FAB_PLL_LOCK(LOCK), .FAB_RXACTIVE(VCC_net_1), 
        .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(GND_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(CORERESETP_0_RESET_N_F2M), 
        .XCLK_FAB(VCC_net_1), .CLK_BASE(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .CLK_MDDR_APB(VCC_net_1), .F_ARADDR_HADDR1({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_ARBURST_HTRANS1({GND_net_1, GND_net_1}), 
        .F_ARID_HSEL1({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_ARLEN_HBURST1({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_ARLOCK_HMASTLOCK1({GND_net_1, GND_net_1}), .F_ARSIZE_HSIZE1({
        GND_net_1, GND_net_1}), .F_ARVALID_HWRITE1(GND_net_1), 
        .F_AWADDR_HADDR0({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_AWBURST_HTRANS0({
        GND_net_1, GND_net_1}), .F_AWID_HSEL0({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_AWLEN_HBURST0({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_AWLOCK_HMASTLOCK0({GND_net_1, 
        GND_net_1}), .F_AWSIZE_HSIZE0({GND_net_1, GND_net_1}), 
        .F_AWVALID_HWRITE0(GND_net_1), .F_BREADY(GND_net_1), 
        .F_RMW_AXI(GND_net_1), .F_RREADY(GND_net_1), .F_WDATA_HWDATA01({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .F_WID_HREADY01({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .F_WLAST(
        GND_net_1), .F_WSTRB({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_WVALID(GND_net_1), .FPGA_MDDR_ARESET_N(VCC_net_1), 
        .MDDR_FABRIC_PADDR({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .MDDR_FABRIC_PENABLE(VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), 
        .MDDR_FABRIC_PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PWRITE(
        VCC_net_1), .PRESET_N(GND_net_1), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), .MGPIO25A_IN(
        GND_net_1), .MGPIO26A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_CTS_MGPIO13B_IN(GND_net_1), .MMUART1_DCD_MGPIO16B_IN(
        GND_net_1), .MMUART1_DSR_MGPIO14B_IN(GND_net_1), 
        .MMUART1_DTR_MGPIO12B_IN(GND_net_1), .MMUART1_RI_MGPIO15B_IN(
        GND_net_1), .MMUART1_RTS_MGPIO11B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), 
        .SPI0_SS4_MGPIO19A_IN(GND_net_1), .SPI0_SS5_MGPIO20A_IN(
        GND_net_1), .SPI0_SS6_MGPIO21A_IN(GND_net_1), 
        .SPI0_SS7_MGPIO22A_IN(GND_net_1), .SPI1_SCK_IN(GND_net_1), 
        .SPI1_SDI_MGPIO11A_IN(GND_net_1), .SPI1_SDO_MGPIO12A_IN(
        GND_net_1), .SPI1_SS0_MGPIO13A_IN(GND_net_1), 
        .SPI1_SS1_MGPIO14A_IN(GND_net_1), .SPI1_SS2_MGPIO15A_IN(
        GND_net_1), .SPI1_SS3_MGPIO16A_IN(GND_net_1), 
        .SPI1_SS4_MGPIO17A_IN(GND_net_1), .SPI1_SS5_MGPIO18A_IN(
        GND_net_1), .SPI1_SS6_MGPIO23A_IN(GND_net_1), 
        .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(GND_net_1), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc274, nc275, 
        nc276, nc277, nc278, nc279, nc280, nc281, nc282, nc283, nc284, 
        nc285, nc286, nc287, nc288, nc289}), .DRAM_BA({nc290, nc291, 
        nc292}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc293, nc294, nc295}), .DRAM_DQ_OUT({nc296, 
        nc297, nc298, nc299, nc300, nc301, nc302, nc303, nc304, nc305, 
        nc306, nc307, nc308, nc309, nc310, nc311, nc312, nc313}), 
        .DRAM_DQS_OUT({nc314, nc315, nc316}), .DRAM_FIFO_WE_OUT({nc317, 
        nc318}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), .MGPIO25A_OUT(), 
        .MGPIO26A_OUT(), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_CTS_MGPIO13B_OUT(), .MMUART1_DCD_MGPIO16B_OUT(), 
        .MMUART1_DSR_MGPIO14B_OUT(), .MMUART1_DTR_MGPIO12B_OUT(), 
        .MMUART1_RI_MGPIO15B_OUT(), .MMUART1_RTS_MGPIO11B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI0_SS4_MGPIO19A_OUT(), 
        .SPI0_SS5_MGPIO20A_OUT(), .SPI0_SS6_MGPIO21A_OUT(), 
        .SPI0_SS7_MGPIO22A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc319, nc320, 
        nc321}), .DRAM_DQ_OE({nc322, nc323, nc324, nc325, nc326, nc327, 
        nc328, nc329, nc330, nc331, nc332, nc333, nc334, nc335, nc336, 
        nc337, nc338, nc339}), .DRAM_DQS_OE({nc340, nc341, nc342}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), .MGPIO25A_OE(), 
        .MGPIO26A_OE(), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), .MMUART1_CTS_MGPIO13B_OE()
        , .MMUART1_DCD_MGPIO16B_OE(), .MMUART1_DSR_MGPIO14B_OE(), 
        .MMUART1_DTR_MGPIO12B_OE(), .MMUART1_RI_MGPIO15B_OE(), 
        .MMUART1_RTS_MGPIO11B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI0_SS4_MGPIO19A_OE(), 
        .SPI0_SS5_MGPIO20A_OE(), .SPI0_SS6_MGPIO21A_OE(), 
        .SPI0_SS7_MGPIO22A_OE(), .SPI1_SCK_OE(), .SPI1_SDI_MGPIO11A_OE(
        ), .SPI1_SDO_MGPIO12A_OE(), .SPI1_SS0_MGPIO13A_OE(), 
        .SPI1_SS1_MGPIO14A_OE(), .SPI1_SS2_MGPIO15A_OE(), 
        .SPI1_SS3_MGPIO16A_OE(), .SPI1_SS4_MGPIO17A_OE(), 
        .SPI1_SS5_MGPIO18A_OE(), .SPI1_SS6_MGPIO23A_OE(), 
        .SPI1_SS7_MGPIO24A_OE(), .USBC_XCLK_OE());
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_23 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[24] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[24]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_1 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[2] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[2]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_22 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[23] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[23]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_20 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[21] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[21]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_25 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[26] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[26]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_5 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[6] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[6]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_7 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[8] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[8]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_6 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[7] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[7]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_30 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[31] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[31]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_2 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[3] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[3]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_8 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[9] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[9]));
    CFG3 #( .INIT(8'h40) )  MSS_ADLIB_INST_RNII8IJ_17 (.A(N_546), .B(
        \CoreAHBLite_0_AHBmslave16_HRDATA[18] ), .C(m0s16DataSel), .Y(
        AHB_IF_0_BIF_1_HRDATA[18]));
    
endmodule


module eSRAM_eNVM_access(
       AHB_IF_0_BIF_1_HADDR,
       AHB_IF_0_BIF_1_HTRANS,
       AHB_IF_0_BIF_1_HWDATA,
       AHB_IF_0_BIF_1_HRDATA,
       DEVRST_N,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       eSRAM_eNVM_access_0_HPMS_READY,
       AHB_IF_0_BIF_1_HWRITE,
       defSlaveSMCurrentState,
       defSlaveSMNextState,
       N_53,
       N_546,
       HREADY_M_0_iv_i_0,
       FAB_RESET_N_c
    );
input  [31:2] AHB_IF_0_BIF_1_HADDR;
input  [1:1] AHB_IF_0_BIF_1_HTRANS;
input  [31:0] AHB_IF_0_BIF_1_HWDATA;
output [31:0] AHB_IF_0_BIF_1_HRDATA;
input  DEVRST_N;
output eSRAM_eNVM_access_0_FIC_0_CLK;
output eSRAM_eNVM_access_0_HPMS_READY;
input  AHB_IF_0_BIF_1_HWRITE;
output defSlaveSMCurrentState;
output defSlaveSMNextState;
output N_53;
output N_546;
output HREADY_M_0_iv_i_0;
input  FAB_RESET_N_c;

    wire SYSRESET_POR_net_1, LOCK, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \sdec_raw_2[0] , \CoreAHBLite_0_AHBmslave16_HWDATA[0] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , m0s16DataSel, N_60, 
        g0_1, CoreAHBLite_0_AHBmslave16_HREADY, N_260, N_33_i_0, 
        N_108_i_0, N_118_i_0, N_116_i_0, N_114_i_0, N_112_i_0, 
        N_110_i_0, N_39_i_0, N_37_i_0, N_106_i_0, N_104_i_0, N_102_i_0, 
        N_100_i_0, N_98_i_0, N_96_i_0, N_94_i_0, N_92_i_0, N_90_i_0, 
        N_88_i_0, N_86_i_0, N_17_i_0, N_16_i_0, N_15_i_0, N_78_i_0, 
        N_14_i_0, N_74_i_0, N_72_i_0, N_70_i_0, N_68_i_0, N_13_i_0, 
        N_64_i_0, N_12_i_0, N_11_i_0, 
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CORERESETP_0_RESET_N_F2M, 
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F, GND_net_1, 
        VCC_net_1;
    
    eSRAM_eNVM_access_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    CoreResetP_Z6_layer0 CORERESETP_0 (.eSRAM_eNVM_access_0_HPMS_READY(
        eSRAM_eNVM_access_0_HPMS_READY), 
        .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N(
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .FAB_RESET_N_c(FAB_RESET_N_c), .CORERESETP_0_RESET_N_F2M(
        CORERESETP_0_RESET_N_F2M), .SYSRESET_POR(SYSRESET_POR_net_1), 
        .eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F(
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F));
    CoreAHBLite_Z5_layer0 CoreAHBLite_0 (.AHB_IF_0_BIF_1_HADDR({
        AHB_IF_0_BIF_1_HADDR[31], AHB_IF_0_BIF_1_HADDR[30], 
        AHB_IF_0_BIF_1_HADDR[29], AHB_IF_0_BIF_1_HADDR[28], 
        AHB_IF_0_BIF_1_HADDR[27], AHB_IF_0_BIF_1_HADDR[26], 
        AHB_IF_0_BIF_1_HADDR[25], AHB_IF_0_BIF_1_HADDR[24], 
        AHB_IF_0_BIF_1_HADDR[23], AHB_IF_0_BIF_1_HADDR[22], 
        AHB_IF_0_BIF_1_HADDR[21], AHB_IF_0_BIF_1_HADDR[20], 
        AHB_IF_0_BIF_1_HADDR[19], AHB_IF_0_BIF_1_HADDR[18], 
        AHB_IF_0_BIF_1_HADDR[17], AHB_IF_0_BIF_1_HADDR[16], 
        AHB_IF_0_BIF_1_HADDR[15], AHB_IF_0_BIF_1_HADDR[14], 
        AHB_IF_0_BIF_1_HADDR[13], AHB_IF_0_BIF_1_HADDR[12], 
        AHB_IF_0_BIF_1_HADDR[11], AHB_IF_0_BIF_1_HADDR[10], 
        AHB_IF_0_BIF_1_HADDR[9], AHB_IF_0_BIF_1_HADDR[8], 
        AHB_IF_0_BIF_1_HADDR[7], AHB_IF_0_BIF_1_HADDR[6], 
        AHB_IF_0_BIF_1_HADDR[5], AHB_IF_0_BIF_1_HADDR[4], 
        AHB_IF_0_BIF_1_HADDR[3], AHB_IF_0_BIF_1_HADDR[2]}), 
        .AHB_IF_0_BIF_1_HTRANS({AHB_IF_0_BIF_1_HTRANS[1]}), 
        .sdec_raw_2({\sdec_raw_2[0] }), .AHB_IF_0_BIF_1_HWDATA({
        AHB_IF_0_BIF_1_HWDATA[31], AHB_IF_0_BIF_1_HWDATA[30], 
        AHB_IF_0_BIF_1_HWDATA[29], AHB_IF_0_BIF_1_HWDATA[28], 
        AHB_IF_0_BIF_1_HWDATA[27], AHB_IF_0_BIF_1_HWDATA[26], 
        AHB_IF_0_BIF_1_HWDATA[25], AHB_IF_0_BIF_1_HWDATA[24], 
        AHB_IF_0_BIF_1_HWDATA[23], AHB_IF_0_BIF_1_HWDATA[22], 
        AHB_IF_0_BIF_1_HWDATA[21], AHB_IF_0_BIF_1_HWDATA[20], 
        AHB_IF_0_BIF_1_HWDATA[19], AHB_IF_0_BIF_1_HWDATA[18], 
        AHB_IF_0_BIF_1_HWDATA[17], AHB_IF_0_BIF_1_HWDATA[16], 
        AHB_IF_0_BIF_1_HWDATA[15], AHB_IF_0_BIF_1_HWDATA[14], 
        AHB_IF_0_BIF_1_HWDATA[13], AHB_IF_0_BIF_1_HWDATA[12], 
        AHB_IF_0_BIF_1_HWDATA[11], AHB_IF_0_BIF_1_HWDATA[10], 
        AHB_IF_0_BIF_1_HWDATA[9], AHB_IF_0_BIF_1_HWDATA[8], 
        AHB_IF_0_BIF_1_HWDATA[7], AHB_IF_0_BIF_1_HWDATA[6], 
        AHB_IF_0_BIF_1_HWDATA[5], AHB_IF_0_BIF_1_HWDATA[4], 
        AHB_IF_0_BIF_1_HWDATA[3], AHB_IF_0_BIF_1_HWDATA[2], 
        AHB_IF_0_BIF_1_HWDATA[1], AHB_IF_0_BIF_1_HWDATA[0]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[0] }), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .m0s16DataSel(m0s16DataSel), .AHB_IF_0_BIF_1_HWRITE(
        AHB_IF_0_BIF_1_HWRITE), .N_60(N_60), .defSlaveSMCurrentState(
        defSlaveSMCurrentState), .defSlaveSMNextState(
        defSlaveSMNextState), .g0_1(g0_1), .N_53(N_53), .N_546(N_546), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .HREADY_M_0_iv_i_0(
        HREADY_M_0_iv_i_0), .N_260(N_260), .N_33_i_0(N_33_i_0), 
        .N_108_i_0(N_108_i_0), .N_118_i_0(N_118_i_0), .N_116_i_0(
        N_116_i_0), .N_114_i_0(N_114_i_0), .N_112_i_0(N_112_i_0), 
        .N_110_i_0(N_110_i_0), .N_39_i_0(N_39_i_0), .N_37_i_0(N_37_i_0)
        , .N_106_i_0(N_106_i_0), .N_104_i_0(N_104_i_0), .N_102_i_0(
        N_102_i_0), .N_100_i_0(N_100_i_0), .N_98_i_0(N_98_i_0), 
        .N_96_i_0(N_96_i_0), .N_94_i_0(N_94_i_0), .N_92_i_0(N_92_i_0), 
        .N_90_i_0(N_90_i_0), .N_88_i_0(N_88_i_0), .N_86_i_0(N_86_i_0), 
        .N_17_i_0(N_17_i_0), .N_16_i_0(N_16_i_0), .N_15_i_0(N_15_i_0), 
        .N_78_i_0(N_78_i_0), .N_14_i_0(N_14_i_0), .N_74_i_0(N_74_i_0), 
        .N_72_i_0(N_72_i_0), .N_70_i_0(N_70_i_0), .N_68_i_0(N_68_i_0), 
        .N_13_i_0(N_13_i_0), .N_64_i_0(N_64_i_0), .N_12_i_0(N_12_i_0), 
        .N_11_i_0(N_11_i_0));
    VCC VCC (.Y(VCC_net_1));
    eSRAM_eNVM_access_CCC_0_FCCC CCC_0 (.eSRAM_eNVM_access_0_FIC_0_CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .LOCK(LOCK), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    GND GND (.Y(GND_net_1));
    eSRAM_eNVM_access_HPMS eSRAM_eNVM_access_HPMS_0 (.sdec_raw_2({
        \sdec_raw_2[0] }), .AHB_IF_0_BIF_1_HRDATA({
        AHB_IF_0_BIF_1_HRDATA[31], AHB_IF_0_BIF_1_HRDATA[30], 
        AHB_IF_0_BIF_1_HRDATA[29], AHB_IF_0_BIF_1_HRDATA[28], 
        AHB_IF_0_BIF_1_HRDATA[27], AHB_IF_0_BIF_1_HRDATA[26], 
        AHB_IF_0_BIF_1_HRDATA[25], AHB_IF_0_BIF_1_HRDATA[24], 
        AHB_IF_0_BIF_1_HRDATA[23], AHB_IF_0_BIF_1_HRDATA[22], 
        AHB_IF_0_BIF_1_HRDATA[21], AHB_IF_0_BIF_1_HRDATA[20], 
        AHB_IF_0_BIF_1_HRDATA[19], AHB_IF_0_BIF_1_HRDATA[18], 
        AHB_IF_0_BIF_1_HRDATA[17], AHB_IF_0_BIF_1_HRDATA[16], 
        AHB_IF_0_BIF_1_HRDATA[15], AHB_IF_0_BIF_1_HRDATA[14], 
        AHB_IF_0_BIF_1_HRDATA[13], AHB_IF_0_BIF_1_HRDATA[12], 
        AHB_IF_0_BIF_1_HRDATA[11], AHB_IF_0_BIF_1_HRDATA[10], 
        AHB_IF_0_BIF_1_HRDATA[9], AHB_IF_0_BIF_1_HRDATA[8], 
        AHB_IF_0_BIF_1_HRDATA[7], AHB_IF_0_BIF_1_HRDATA[6], 
        AHB_IF_0_BIF_1_HRDATA[5], AHB_IF_0_BIF_1_HRDATA[4], 
        AHB_IF_0_BIF_1_HRDATA[3], AHB_IF_0_BIF_1_HRDATA[2], 
        AHB_IF_0_BIF_1_HRDATA[1], AHB_IF_0_BIF_1_HRDATA[0]}), 
        .CoreAHBLite_0_AHBmslave16_HWDATA({
        \CoreAHBLite_0_AHBmslave16_HWDATA[31] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[30] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[29] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[28] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[27] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[26] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[25] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[24] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[23] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[22] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[21] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[20] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[19] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[18] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[17] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[16] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[15] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[14] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[13] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[12] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[11] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[10] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[9] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[8] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[7] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[6] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[5] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[4] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[3] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[2] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[1] , 
        \CoreAHBLite_0_AHBmslave16_HWDATA[0] }), .N_60(N_60), 
        .CoreAHBLite_0_AHBmslave16_HREADY(
        CoreAHBLite_0_AHBmslave16_HREADY), .g0_1(g0_1), .N_546(N_546), 
        .m0s16DataSel(m0s16DataSel), 
        .eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N(
        eSRAM_eNVM_access_HPMS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F(
        eSRAM_eNVM_access_HPMS_TMP_0_MSS_RESET_N_M2F), .N_11_i_0(
        N_11_i_0), .N_12_i_0(N_12_i_0), .N_64_i_0(N_64_i_0), .N_13_i_0(
        N_13_i_0), .N_68_i_0(N_68_i_0), .N_70_i_0(N_70_i_0), .N_72_i_0(
        N_72_i_0), .N_74_i_0(N_74_i_0), .N_14_i_0(N_14_i_0), .N_78_i_0(
        N_78_i_0), .N_15_i_0(N_15_i_0), .N_16_i_0(N_16_i_0), .N_17_i_0(
        N_17_i_0), .N_86_i_0(N_86_i_0), .N_88_i_0(N_88_i_0), .N_90_i_0(
        N_90_i_0), .N_92_i_0(N_92_i_0), .N_94_i_0(N_94_i_0), .N_96_i_0(
        N_96_i_0), .N_98_i_0(N_98_i_0), .N_100_i_0(N_100_i_0), 
        .N_102_i_0(N_102_i_0), .N_104_i_0(N_104_i_0), .N_106_i_0(
        N_106_i_0), .N_37_i_0(N_37_i_0), .N_39_i_0(N_39_i_0), 
        .N_108_i_0(N_108_i_0), .N_110_i_0(N_110_i_0), .N_112_i_0(
        N_112_i_0), .N_114_i_0(N_114_i_0), .N_260(N_260), .N_116_i_0(
        N_116_i_0), .N_33_i_0(N_33_i_0), .N_118_i_0(N_118_i_0), .LOCK(
        LOCK), .CORERESETP_0_RESET_N_F2M(CORERESETP_0_RESET_N_F2M), 
        .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    
endmodule


module eSRAM_eNVM_RW(
       eSRAM_eNVM_RW_0_ram_waddr,
       eSRAM_eNVM_RW_0_ram_wdata,
       AHB_IF_0_DATAOUT,
       state,
       eSRAM_eNVM_RW_0_ADDR,
       eSRAM_eNVM_RW_0_DATAOUT,
       eSRAM_eNVM_access_0_HPMS_READY,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       eSRAM_eNVM_RW_0_WRITE,
       eSRAM_eNVM_RW_0_READ,
       eSRAM_eNVM_RW_0_ram_wen,
       start_esram_c,
       AHB_IF_0_AHB_BUSY,
       AHB_IF_0_VALID
    );
output [4:0] eSRAM_eNVM_RW_0_ram_waddr;
output [31:0] eSRAM_eNVM_RW_0_ram_wdata;
input  [31:0] AHB_IF_0_DATAOUT;
input  [0:0] state;
output [31:2] eSRAM_eNVM_RW_0_ADDR;
output [31:0] eSRAM_eNVM_RW_0_DATAOUT;
input  eSRAM_eNVM_access_0_HPMS_READY;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
output eSRAM_eNVM_RW_0_WRITE;
output eSRAM_eNVM_RW_0_READ;
output eSRAM_eNVM_RW_0_ram_wen;
input  start_esram_c;
input  AHB_IF_0_AHB_BUSY;
input  AHB_IF_0_VALID;

    wire VCC_net_1, N_374_i_0, ram_waddre, GND_net_1, N_376_i_0, 
        N_372_i_0, N_373_i_0, \data_cnt[3]_net_1 , N_322_i_0, 
        \current_state_RNI6JBF1[6]_net_1 , \data_cnt[4]_net_1 , 
        N_323_i_0, N_9_i_0, \data_cnt[0]_net_1 , N_453, 
        \data_cnt[1]_net_1 , N_320_i_0, \data_cnt[2]_net_1 , N_321_i_0, 
        N_149_i_0, N_793_i_0, N_393_i_0, N_379_i_0, N_391_i_0, 
        envm_release_reg_net_1, \current_state[9]_net_1 , 
        un40_0_0_0_net_1, N_292, N_388_i_0, \current_state[6]_net_1 , 
        N_331_i_0, \current_state[7]_net_1 , \current_state_ns[7] , 
        \current_state[8]_net_1 , \current_state_ns[8] , 
        \current_state_ns[9] , \data_13[31] , \current_state_ns[10] , 
        \current_state[11]_net_1 , N_337_i_0, 
        \current_state[12]_net_1 , \current_state_ns[12] , 
        \current_state[13]_net_1 , N_340_i_0, 
        \current_state[14]_net_1 , N_342_i_0, 
        \current_state[15]_net_1 , \current_state_ns[15] , 
        \current_state[16]_net_1 , \current_state_ns[16] , 
        \current_state[0]_net_1 , \current_state_ns[0] , 
        \current_state[1]_net_1 , \current_state_ns_i_i_0[1]_net_1 , 
        \current_state[2]_net_1 , \current_state_ns[2] , 
        \current_state[3]_net_1 , \current_state_ns[3] , 
        \current_state[4]_net_1 , \current_state_ns_i_i_0[4]_net_1 , 
        \current_state[5]_net_1 , \current_state_ns[5] , 
        start_esram_reg_net_1, start_envm_reg1_net_1, 
        start_esram_reg1_net_1, start_envm_reg2_net_1, 
        start_esram_reg2_net_1, \addr_temp_lm[2] , N_40, 
        \addr_temp_lm[3] , \addr_temp_lm[4] , \addr_temp_lm[5] , 
        \addr_temp_lm[6] , \addr_temp_lm[7] , \addr_temp_lm[8] , 
        \addr_temp_lm[9] , \addr_temp_lm[10] , \addr_temp_lm[11] , 
        \addr_temp_lm[12] , \addr_temp_lm[13] , \addr_temp_lm[14] , 
        \addr_temp_lm[15] , \addr_temp_lm[16] , \addr_temp_lm[17] , 
        \addr_temp_lm[18] , \addr_temp_lm[19] , \addr_temp_lm[20] , 
        \addr_temp_lm[21] , \addr_temp_lm[22] , \addr_temp_lm[23] , 
        \addr_temp_lm[24] , \addr_temp_lm[25] , \addr_temp_lm[26] , 
        \addr_temp_lm[27] , \addr_temp_lm[28] , \addr_temp_lm[29] , 
        \addr_temp_lm[30] , \addr_temp_lm[31] , \data_lm[0] , 
        N_141_i_0, \data_lm[1] , \data_lm[2] , \data_lm[3] , 
        \data_lm[4] , \data_lm[5] , \data_lm[6] , \data_lm[7] , 
        \data_lm[8] , \data_lm[9] , \data_lm[10] , \data_lm[11] , 
        \data_lm[12] , \data_lm[13] , \data_lm[14] , \data_lm[15] , 
        \data_lm[16] , \data_lm[17] , \data_lm[18] , \data_lm[19] , 
        \data_lm[20] , \data_lm[21] , \data_lm[22] , \data_lm[23] , 
        \data_lm[24] , \data_lm[25] , \data_lm[26] , \data_lm[27] , 
        \data_lm[28] , \data_lm[29] , \data_lm[30] , \data_lm[31] , 
        data_s_71_FCO, \data_cry[1]_net_1 , \data_s[1] , 
        \data_cry[2]_net_1 , \data_s[2] , \data_cry[3]_net_1 , 
        \data_s[3] , \data_cry[4]_net_1 , \data_s[4] , 
        \data_cry[5]_net_1 , \data_s[5] , \data_cry[6]_net_1 , 
        \data_s[6] , \data_cry[7]_net_1 , \data_s[7] , 
        \data_cry[8]_net_1 , \data_s[8] , \data_cry[9]_net_1 , 
        \data_s[9] , \data_cry[10]_net_1 , \data_s[10] , 
        \data_cry[11]_net_1 , \data_s[11] , \data_cry[12]_net_1 , 
        \data_s[12] , \data_cry[13]_net_1 , \data_s[13] , 
        \data_cry[14]_net_1 , \data_s[14] , \data_cry[15]_net_1 , 
        \data_s[15] , \data_cry[16]_net_1 , \data_s[16] , 
        \data_cry[17]_net_1 , \data_s[17] , \data_cry[18]_net_1 , 
        \data_s[18] , \data_cry[19]_net_1 , \data_s[19] , 
        \data_cry[20]_net_1 , \data_s[20] , \data_cry[21]_net_1 , 
        \data_s[21] , \data_cry[22]_net_1 , \data_s[22] , 
        \data_cry[23]_net_1 , \data_s[23] , \data_cry[24]_net_1 , 
        \data_s[24] , \data_cry[25]_net_1 , \data_s[25] , 
        \data_cry[26]_net_1 , \data_s[26] , \data_cry[27]_net_1 , 
        \data_s[27] , \data_cry[28]_net_1 , \data_s[28] , 
        \data_cry[29]_net_1 , \data_s[29] , \data_s[31]_net_1 , 
        \data_cry[30]_net_1 , \data_s[30] , addr_temp_s_72_FCO, 
        \addr_temp_cry[3]_net_1 , \addr_temp_s[3] , 
        \addr_temp_cry[4]_net_1 , \addr_temp_s[4] , 
        \addr_temp_cry[5]_net_1 , \addr_temp_s[5] , 
        \addr_temp_cry[6]_net_1 , \addr_temp_s[6] , 
        \addr_temp_cry[7]_net_1 , \addr_temp_s[7] , 
        \addr_temp_cry[8]_net_1 , \addr_temp_s[8] , 
        \addr_temp_cry[9]_net_1 , \addr_temp_s[9] , 
        \addr_temp_cry[10]_net_1 , \addr_temp_s[10] , 
        \addr_temp_cry[11]_net_1 , \addr_temp_s[11] , 
        \addr_temp_cry[12]_net_1 , \addr_temp_s[12] , 
        \addr_temp_cry[13]_net_1 , \addr_temp_s[13] , 
        \addr_temp_cry[14]_net_1 , \addr_temp_s[14] , 
        \addr_temp_cry[15]_net_1 , \addr_temp_s[15] , 
        \addr_temp_cry[16]_net_1 , \addr_temp_s[16] , 
        \addr_temp_cry[17]_net_1 , \addr_temp_s[17] , 
        \addr_temp_cry[18]_net_1 , \addr_temp_s[18] , 
        \addr_temp_cry[19]_net_1 , \addr_temp_s[19] , 
        \addr_temp_cry[20]_net_1 , \addr_temp_s[20] , 
        \addr_temp_cry[21]_net_1 , \addr_temp_s[21] , 
        \addr_temp_cry[22]_net_1 , \addr_temp_s[22] , 
        \addr_temp_cry[23]_net_1 , \addr_temp_s[23] , 
        \addr_temp_cry[24]_net_1 , \addr_temp_s[24] , 
        \addr_temp_cry[25]_net_1 , \addr_temp_s[25] , 
        \addr_temp_cry[26]_net_1 , \addr_temp_s[26] , 
        \addr_temp_cry[27]_net_1 , \addr_temp_s[27] , 
        \addr_temp_cry[28]_net_1 , \addr_temp_s[28] , 
        \addr_temp_cry[29]_net_1 , \addr_temp_s[29] , 
        \addr_temp_s[31]_net_1 , \addr_temp_cry[30]_net_1 , 
        \addr_temp_s[30] , \data_13[6] , N_337, N_387, N_341, 
        un1_addr_temp_8_sqmuxa_2_i_i_i_1, N_340, N_349, N_272, N_357, 
        N_822, \addr_temp_lm_0_1_0[2]_net_1 , 
        \addr_temp_lm_0_1[7]_net_1 , N_448, N_393_i_1, N_409, N_531, 
        N_532, N_407_2, \data_lm_0_1_0[0]_net_1 , 
        \current_state_RNIHJVS3[2]_net_1 , N_333, 
        un1_current_state_20_i_0_0_a2_0_2_net_1, 
        un1_current_state_20_i_0_0_a2_0_4_net_1, 
        \addr_temp_cnst_i_a2_0_i_a2_0_0[8]_net_1 , N_379, 
        un1_current_state_20_i_0_0_a2_0_0_net_1, 
        un1_current_state_16_0_0_i_0_0_a2_1_0, 
        un1_current_state_13_i_0_0_a2_0_net_1, 
        ram_wdata_0_sqmuxa_i_a6_0_4_0_net_1, esram_select_net_1, N_339, 
        N_355, N_343, N_513, ram_wdata_0_sqmuxa_i_0_net_1, 
        ram_wdata_0_sqmuxa_i_a6_1_3_net_1, un1_READ6_3_0_0_0_2, 
        un1_current_state_16_0_0_i_0_0_a2_0_0, N_370_i_i_0_a2_1_2, 
        \addr_temp_cnst_i_a2_0_i_o2_1_0[8]_net_1 , 
        un1_READ_1_sqmuxa_2_i_0_a3_2_net_1, 
        un1_READ_1_sqmuxa_2_i_0_a3_1_net_1, 
        ram_wdata_0_sqmuxa_i_a6_3_2_net_1, 
        ram_wdata_0_sqmuxa_i_a6_0_4_2_net_1, 
        un1_current_state_16_0_0_i_0_0_a2_2_0, 
        un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3_net_1, 
        un1_READ_1_sqmuxa_2_i_0_a3_2_2_net_1, 
        \addr_temp_cnst_0_a2_i_0_o2_a0[19]_net_1 , 
        un1_addr_temp_8_sqmuxa_2_i_i_o2_3_0_c, N_439, N_498, N_499, 
        N_511, N_360, N_516, N_314, N_352, 
        ram_wdata_0_sqmuxa_i_a6_1_4_net_1, 
        un1_current_state_16_0_0_i_0_0_a2_1_2, N_370_i_i_0_a2_1_3, 
        \current_state_ns_i_0_0_0[13]_net_1 , 
        ram_wdata_0_sqmuxa_i_a6_3_net_1, N_465, N_461, N_103, N_335, 
        \addr_temp_cnst_0_a2_i_a6_0[30]_net_1 , N_362, N_241, 
        un1_current_state_16_0_0_i_0_0_0, N_512, N_384, 
        ram_wdata_0_sqmuxa_i_2_tz_net_1, 
        un1_READ_1_sqmuxa_2_i_0_0_net_1, N_530, N_410, N_347_i, N_514, 
        \data_13[7] , un1_current_state_16_0_0_i_0_0_1, N_370_i_i_0_0, 
        un1_current_state_20_i_0_0_0_net_1;
    
    CFG2 #( .INIT(4'h7) )  ram_waddr_n2_0_o2 (.A(
        eSRAM_eNVM_RW_0_ram_waddr[0]), .B(eSRAM_eNVM_RW_0_ram_waddr[1])
        , .Y(N_343));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[24]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[24]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[23]_net_1 ), .S(\data_s[24] ), .Y(), .FCO(
        \data_cry[24]_net_1 ));
    CFG4 #( .INIT(16'hF888) )  \current_state_ns_0_0[9]  (.A(
        \current_state[8]_net_1 ), .B(AHB_IF_0_DATAOUT[0]), .C(
        \current_state[9]_net_1 ), .D(N_341), .Y(\current_state_ns[9] )
        );
    CFG4 #( .INIT(16'hCA0A) )  \addr_temp_lm_0[4]  (.A(
        \addr_temp_s[4] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_337), .Y(\addr_temp_lm[4] ));
    CFG4 #( .INIT(16'hCAC0) )  \current_state_ns_0_0[7]  (.A(
        \current_state[6]_net_1 ), .B(\current_state[7]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_514), .Y(\current_state_ns[7] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[26]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[26]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[25]_net_1 ), .S(\addr_temp_s[26] ), .Y(), .FCO(
        \addr_temp_cry[26]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[12]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[11]_net_1 ), .S(\addr_temp_s[12] ), .Y(), .FCO(
        \addr_temp_cry[12]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \data_lm_0_1_0[0]  (.A(N_333), .B(
        \current_state[4]_net_1 ), .Y(\data_lm_0_1_0[0]_net_1 ));
    CFG4 #( .INIT(16'hA0CC) )  \addr_temp_lm_0[16]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\addr_temp_s[16] ), .C(
        \data_13[6] ), .D(N_822), .Y(\addr_temp_lm[16] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[20]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[20]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[19]_net_1 ), .S(\addr_temp_s[20] ), .Y(), .FCO(
        \addr_temp_cry[20]_net_1 ));
    SLE \data[5]  (.D(\data_lm[5] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[5]));
    SLE \addr_temp[25]  (.D(\addr_temp_lm[25] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[25]));
    SLE \ram_wdata[9]  (.D(AHB_IF_0_DATAOUT[9]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[9]));
    CFG4 #( .INIT(16'h55C3) )  \ram_waddr_RNO[4]  (.A(
        \current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ram_waddr[4]), 
        .C(N_362), .D(N_384), .Y(N_376_i_0));
    CFG4 #( .INIT(16'h8F80) )  \addr_temp_lm_0[10]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\current_state[9]_net_1 ), 
        .C(N_822), .D(\addr_temp_s[10] ), .Y(\addr_temp_lm[10] ));
    SLE \addr_temp[16]  (.D(\addr_temp_lm[16] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[16]));
    CFG2 #( .INIT(4'h1) )  ram_wdata_0_sqmuxa_i_a6_0_4_0 (.A(
        \current_state[12]_net_1 ), .B(\current_state[6]_net_1 ), .Y(
        ram_wdata_0_sqmuxa_i_a6_0_4_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[29]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[29]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[28]_net_1 ), .S(\data_s[29] ), .Y(), .FCO(
        \data_cry[29]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[28]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[28]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[27]_net_1 ), .S(\data_s[28] ), .Y(), .FCO(
        \data_cry[28]_net_1 ));
    CFG4 #( .INIT(16'hCA0A) )  \addr_temp_lm_0[3]  (.A(
        \addr_temp_s[3] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_387), .Y(\addr_temp_lm[3] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[3]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        addr_temp_s_72_FCO), .S(\addr_temp_s[3] ), .Y(), .FCO(
        \addr_temp_cry[3]_net_1 ));
    SLE \current_state[2]  (.D(\current_state_ns[2] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[2]_net_1 ));
    CFG4 #( .INIT(16'hFFF4) )  \addr_temp_cnst_i_a2_i_0_o2[3]  (.A(
        AHB_IF_0_AHB_BUSY), .B(\current_state[7]_net_1 ), .C(
        \data_13[6] ), .D(N_337), .Y(N_387));
    CFG4 #( .INIT(16'h0007) )  WRITE_RNO (.A(N_514), .B(
        un1_current_state_16_0_0_i_0_0_a2_1_2), .C(N_410), .D(
        un1_current_state_16_0_0_i_0_0_1), .Y(N_793_i_0));
    CFG3 #( .INIT(8'h20) )  un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2 (.A(
        eSRAM_eNVM_RW_0_ram_waddr[2]), .B(eSRAM_eNVM_RW_0_ram_waddr[0])
        , .C(un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3_net_1), .Y(N_103));
    CFG4 #( .INIT(16'hA0CC) )  \addr_temp_lm_0[15]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\addr_temp_s[15] ), .C(
        \data_13[6] ), .D(N_822), .Y(\addr_temp_lm[15] ));
    SLE \ram_wdata[23]  (.D(AHB_IF_0_DATAOUT[23]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[23]));
    SLE \data[9]  (.D(\data_lm[9] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[9]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[27]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[27]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[26]_net_1 ), .S(\addr_temp_s[27] ), .Y(), .FCO(
        \addr_temp_cry[27]_net_1 ));
    SLE \addr_temp[26]  (.D(\addr_temp_lm[26] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[26]));
    SLE \data[10]  (.D(\data_lm[10] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[10]));
    SLE \addr_temp[3]  (.D(\addr_temp_lm[3] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[3]));
    SLE \current_state[6]  (.D(N_331_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[6]_net_1 ));
    SLE \addr_temp[13]  (.D(\addr_temp_lm[13] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[13]));
    SLE \data_cnt[2]  (.D(N_321_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        \current_state_RNI6JBF1[6]_net_1 ), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_cnt[2]_net_1 ));
    SLE \ram_wdata[17]  (.D(AHB_IF_0_DATAOUT[17]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[17]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[24]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[24]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[23]_net_1 ), .S(\addr_temp_s[24] ), .Y(), .FCO(
        \addr_temp_cry[24]_net_1 ));
    SLE \data[13]  (.D(\data_lm[13] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[13]));
    SLE \ram_wdata[8]  (.D(AHB_IF_0_DATAOUT[8]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[8]));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[12]  (.A(N_822), .B(
        \addr_temp_s[12] ), .Y(\addr_temp_lm[12] ));
    CFG4 #( .INIT(16'hCC40) )  \addr_temp_cnst_0_a2_i_a6_0[30]  (.A(
        AHB_IF_0_AHB_BUSY), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        \current_state[12]_net_1 ), .D(\data_13[31] ), .Y(
        \addr_temp_cnst_0_a2_i_a6_0[30]_net_1 ));
    SLE \addr_temp[6]  (.D(\addr_temp_lm[6] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[6]));
    SLE \addr_temp[23]  (.D(\addr_temp_lm[23] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[23]));
    CFG4 #( .INIT(16'hCE8A) )  \current_state_ns_i_i_0[4]  (.A(
        \current_state[3]_net_1 ), .B(\current_state[4]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_360), .Y(
        \current_state_ns_i_i_0[4]_net_1 ));
    CFG3 #( .INIT(8'h72) )  \addr_temp_lm_0[30]  (.A(N_822), .B(
        \addr_temp_cnst_0_a2_i_a6_0[30]_net_1 ), .C(\addr_temp_s[30] ), 
        .Y(\addr_temp_lm[30] ));
    CFG2 #( .INIT(4'h1) )  \addr_temp_lm_0_1_0[2]  (.A(\data_13[6] ), 
        .B(N_337), .Y(\addr_temp_lm_0_1_0[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[16]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[16]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[15]_net_1 ), .S(\addr_temp_s[16] ), .Y(), .FCO(
        \addr_temp_cry[16]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[3]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[3] ), .Y(
        \data_lm[3] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[10]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[9]_net_1 ), .S(\addr_temp_s[10] ), .Y(), .FCO(
        \addr_temp_cry[10]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  ram_wdata_0_sqmuxa_i_a6_3 (.A(
        \current_state[8]_net_1 ), .B(\current_state[11]_net_1 ), .C(
        ram_wdata_0_sqmuxa_i_a6_3_2_net_1), .D(\data_13[31] ), .Y(
        ram_wdata_0_sqmuxa_i_a6_3_net_1));
    SLE \addr_temp[7]  (.D(\addr_temp_lm[7] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[7]));
    CFG2 #( .INIT(4'h4) )  \addr_temp_cnst_0_a2_i_0_a2_0[19]  (.A(
        AHB_IF_0_AHB_BUSY), .B(\current_state[12]_net_1 ), .Y(N_513));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[2]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[2] ), .Y(
        \data_lm[2] ));
    CFG3 #( .INIT(8'h8C) )  \ram_waddr_RNIAKOT[2]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[0]), .B(\current_state[14]_net_1 ), 
        .C(eSRAM_eNVM_RW_0_ram_waddr[2]), .Y(
        un1_addr_temp_8_sqmuxa_2_i_i_o2_3_0_c));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[13]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[13] ), .Y(
        \data_lm[13] ));
    SLE \data[4]  (.D(\data_lm[4] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[4]));
    SLE start_esram_reg1 (.D(start_esram_reg_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        start_esram_reg1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[17]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[17]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[16]_net_1 ), .S(\data_s[17] ), .Y(), .FCO(
        \data_cry[17]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  \data_cnt_RNI841P1[4]  (.A(
        \data_cnt[4]_net_1 ), .B(\data_cnt[3]_net_1 ), .C(
        \data_cnt[2]_net_1 ), .D(N_339), .Y(N_514));
    SLE \data[11]  (.D(\data_lm[11] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[11]));
    CFG4 #( .INIT(16'h0002) )  envm_release_reg_RNIPUH21 (.A(
        \current_state[16]_net_1 ), .B(\current_state[4]_net_1 ), .C(
        envm_release_reg_net_1), .D(\current_state[2]_net_1 ), .Y(
        N_531));
    CFG4 #( .INIT(16'h5051) )  \current_state_ns_i_0_0_0[13]  (.A(
        \current_state[13]_net_1 ), .B(AHB_IF_0_VALID), .C(
        AHB_IF_0_AHB_BUSY), .D(\current_state[12]_net_1 ), .Y(
        \current_state_ns_i_0_0_0[13]_net_1 ));
    CFG2 #( .INIT(4'h7) )  data_cnt_n2_i_o2 (.A(\data_cnt[0]_net_1 ), 
        .B(\data_cnt[1]_net_1 ), .Y(N_339));
    SLE \ram_waddr[4]  (.D(N_376_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(ram_waddre), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_ram_waddr[4]));
    CFG4 #( .INIT(16'hFFFE) )  \addr_temp_cnst_0_a2_i_0_o2_1[19]  (.A(
        \data_13[31] ), .B(\current_state[9]_net_1 ), .C(N_513), .D(
        \addr_temp_cnst_0_a2_i_0_o2_a0[19]_net_1 ), .Y(N_272));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[15]  (.A(\data_s[15] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[15] ));
    CFG3 #( .INIT(8'h20) )  un1_current_state_20_i_0_0_a2_0_4 (.A(
        N_532), .B(N_349), .C(un1_current_state_20_i_0_0_a2_0_2_net_1), 
        .Y(un1_current_state_20_i_0_0_a2_0_4_net_1));
    CFG4 #( .INIT(16'h55C3) )  \ram_waddr_RNO[2]  (.A(
        \current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ram_waddr[2]), 
        .C(N_343), .D(N_384), .Y(N_373_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[9]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[9]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[8]_net_1 ), .S(\data_s[9] ), .Y(), .FCO(
        \data_cry[9]_net_1 ));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[17]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[17]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[16]_net_1 ), .S(\addr_temp_s[17] ), .Y(), .FCO(
        \addr_temp_cry[17]_net_1 ));
    SLE \ram_wdata[4]  (.D(AHB_IF_0_DATAOUT[4]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[4]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[7]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[6]_net_1 ), .S(\addr_temp_s[7] ), .Y(), .FCO(
        \addr_temp_cry[7]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \addr_temp_cnst_0_a2_i_0_o2_a0[19]  (.A(
        \current_state[4]_net_1 ), .B(AHB_IF_0_DATAOUT[0]), .C(
        AHB_IF_0_DATAOUT[2]), .D(AHB_IF_0_DATAOUT[1]), .Y(
        \addr_temp_cnst_0_a2_i_0_o2_a0[19]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[18]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[18] ), .Y(
        \data_lm[18] ));
    CFG4 #( .INIT(16'h0001) )  un1_READ_1_sqmuxa_2_i_0_a3_1 (.A(
        \current_state[1]_net_1 ), .B(\current_state[14]_net_1 ), .C(
        \current_state[13]_net_1 ), .D(\current_state[3]_net_1 ), .Y(
        un1_READ_1_sqmuxa_2_i_0_a3_1_net_1));
    CFG2 #( .INIT(4'h1) )  un1_current_state_19_i_0_0_a2_1 (.A(N_355), 
        .B(\current_state[1]_net_1 ), .Y(N_532));
    CFG4 #( .INIT(16'h0008) )  un1_current_state_19_i_0_0_a2_0 (.A(
        un1_current_state_16_0_0_i_0_0_a2_2_0), .B(N_532), .C(
        \current_state[16]_net_1 ), .D(\data_13[31] ), .Y(N_409));
    CFG4 #( .INIT(16'hF2FA) )  \current_state_ns_0_0[0]  (.A(
        \current_state[16]_net_1 ), .B(envm_release_reg_net_1), .C(
        N_465), .D(AHB_IF_0_AHB_BUSY), .Y(\current_state_ns[0] ));
    CFG4 #( .INIT(16'h0001) )  ram_wdata_0_sqmuxa_i_a6_3_2 (.A(
        \current_state[15]_net_1 ), .B(\current_state[14]_net_1 ), .C(
        \current_state[12]_net_1 ), .D(\current_state[9]_net_1 ), .Y(
        ram_wdata_0_sqmuxa_i_a6_3_2_net_1));
    CFG3 #( .INIT(8'h09) )  \data_cnt_RNO[2]  (.A(\data_cnt[2]_net_1 ), 
        .B(N_339), .C(N_314), .Y(N_321_i_0));
    SLE \data_cnt[4]  (.D(N_323_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        \current_state_RNI6JBF1[6]_net_1 ), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_cnt[4]_net_1 ));
    SLE \current_state[5]  (.D(\current_state_ns[5] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[5]_net_1 ));
    CFG2 #( .INIT(4'h1) )  data_cnt_n0_i_a2 (.A(N_314), .B(
        \data_cnt[0]_net_1 ), .Y(N_453));
    CFG2 #( .INIT(4'hE) )  \current_state_RNIDPOE[12]  (.A(
        \current_state[0]_net_1 ), .B(\current_state[12]_net_1 ), .Y(
        N_355));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[14]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[13]_net_1 ), .S(\addr_temp_s[14] ), .Y(), .FCO(
        \addr_temp_cry[14]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[24]  (.A(N_822), .B(
        \addr_temp_s[24] ), .Y(\addr_temp_lm[24] ));
    CFG4 #( .INIT(16'hFFCE) )  \addr_temp_cnst_i_a2_0_i_o2_1[8]  (.A(
        \addr_temp_cnst_i_a2_0_i_a2_0_0[8]_net_1 ), .B(N_337), .C(
        AHB_IF_0_AHB_BUSY), .D(
        \addr_temp_cnst_i_a2_0_i_o2_1_0[8]_net_1 ), .Y(N_357));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[9]  (.A(N_822), .B(
        \addr_temp_s[9] ), .Y(\addr_temp_lm[9] ));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[23]  (.A(\data_s[23] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[23] ));
    CFG4 #( .INIT(16'h0A0E) )  \current_state_RNO[14]  (.A(
        \current_state[14]_net_1 ), .B(\current_state[13]_net_1 ), .C(
        N_103), .D(N_341), .Y(N_342_i_0));
    SLE \data_cnt[1]  (.D(N_320_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        \current_state_RNI6JBF1[6]_net_1 ), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_cnt[1]_net_1 ));
    SLE \ram_wdata[11]  (.D(AHB_IF_0_DATAOUT[11]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[11]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[16]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[16]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[15]_net_1 ), .S(\data_s[16] ), .Y(), .FCO(
        \data_cry[16]_net_1 ));
    SLE \data[24]  (.D(\data_lm[24] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[24]));
    CFG3 #( .INIT(8'h04) )  \current_state_RNI3CDV[2]  (.A(
        \current_state[4]_net_1 ), .B(AHB_IF_0_AHB_BUSY), .C(
        \current_state[2]_net_1 ), .Y(
        un1_current_state_16_0_0_i_0_0_a2_2_0));
    CFG4 #( .INIT(16'h0155) )  READ_RNO_0 (.A(
        un1_current_state_20_i_0_0_0_net_1), .B(N_512), .C(N_511), .D(
        un1_current_state_20_i_0_0_a2_0_4_net_1), .Y(N_391_i_0));
    SLE \ram_wdata[31]  (.D(AHB_IF_0_DATAOUT[31]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[31]));
    SLE \addr_temp[30]  (.D(\addr_temp_lm[30] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[30]));
    ARI1 #( .INIT(20'h4AA00) )  addr_temp_s_72 (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(addr_temp_s_72_FCO));
    CFG4 #( .INIT(16'h0001) )  un1_READ_1_sqmuxa_2_i_0_a3_2_2 (.A(
        AHB_IF_0_VALID), .B(\current_state[3]_net_1 ), .C(
        \current_state[8]_net_1 ), .D(\current_state[12]_net_1 ), .Y(
        un1_READ_1_sqmuxa_2_i_0_a3_2_2_net_1));
    SLE \data[30]  (.D(\data_lm[30] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[30]));
    CFG3 #( .INIT(8'hE0) )  un1_current_state_20_i_0_0_a2 (.A(
        \current_state[8]_net_1 ), .B(\current_state[4]_net_1 ), .C(
        AHB_IF_0_DATAOUT[0]), .Y(N_448));
    SLE \ram_wdata[6]  (.D(AHB_IF_0_DATAOUT[6]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[6]));
    CFG4 #( .INIT(16'hFF40) )  ram_wdata_0_sqmuxa_i_2_tz (.A(
        \current_state[4]_net_1 ), .B(
        ram_wdata_0_sqmuxa_i_a6_0_4_0_net_1), .C(
        ram_wdata_0_sqmuxa_i_a6_0_4_2_net_1), .D(
        ram_wdata_0_sqmuxa_i_a6_3_net_1), .Y(
        ram_wdata_0_sqmuxa_i_2_tz_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[10]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[10]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[9]_net_1 ), .S(\data_s[10] ), .Y(), .FCO(
        \data_cry[10]_net_1 ));
    CFG4 #( .INIT(16'hCACE) )  \current_state_ns_0_0[2]  (.A(
        \current_state[1]_net_1 ), .B(\current_state[2]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(AHB_IF_0_DATAOUT[0]), .Y(
        \current_state_ns[2] ));
    SLE start_esram_reg2 (.D(start_esram_reg1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        start_esram_reg2_net_1));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[30]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[30] ), .Y(
        \data_lm[30] ));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[25]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[25] ), .Y(
        \data_lm[25] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[27]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[27]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[26]_net_1 ), .S(\data_s[27] ), .Y(), .FCO(
        \data_cry[27]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[6]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[6]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[5]_net_1 ), .S(\data_s[6] ), .Y(), .FCO(
        \data_cry[6]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \current_state_RNIH70A1[5]  (.A(
        \current_state[0]_net_1 ), .B(\data_13[31] ), .C(
        \current_state[5]_net_1 ), .D(\current_state[7]_net_1 ), .Y(
        un1_READ6_3_0_0_0_2));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[28]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[28] ), .Y(
        \data_lm[28] ));
    CFG4 #( .INIT(16'h353A) )  \ram_waddr_RNO[1]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[1]), .B(\current_state[0]_net_1 ), 
        .C(N_384), .D(eSRAM_eNVM_RW_0_ram_waddr[0]), .Y(N_372_i_0));
    CFG4 #( .INIT(16'hF5C5) )  \ram_waddr_RNO[0]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[0]), .B(\current_state[12]_net_1 ), 
        .C(N_384), .D(\current_state[9]_net_1 ), .Y(N_9_i_0));
    SLE \data[1]  (.D(\data_lm[1] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[1]));
    CFG2 #( .INIT(4'h1) )  WRITE_RNO_5 (.A(\current_state[5]_net_1 ), 
        .B(\current_state[11]_net_1 ), .Y(
        un1_current_state_16_0_0_i_0_0_a2_1_0));
    CFG3 #( .INIT(8'hAC) )  \data_lm_0[10]  (.A(\data_13[7] ), .B(
        \data_s[10] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[10] ));
    SLE \current_state[16]  (.D(\current_state_ns[16] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[16]_net_1 ));
    SLE \data[6]  (.D(\data_lm[6] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[6]));
    SLE \addr_temp[31]  (.D(\addr_temp_lm[31] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[31]));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[17]  (.A(\data_s[17] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[17] ));
    SLE \data[25]  (.D(\data_lm[25] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[25]));
    CFG3 #( .INIT(8'hEC) )  \current_state_ns_0_0[5]  (.A(
        AHB_IF_0_AHB_BUSY), .B(\data_13[6] ), .C(
        \current_state[5]_net_1 ), .Y(\current_state_ns[5] ));
    SLE \ram_wdata[5]  (.D(AHB_IF_0_DATAOUT[5]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[5]));
    CFG4 #( .INIT(16'h000B) )  
        \addr_temp_cnst_0_a2_i_0_o2_1_RNI42HI1[19]  (.A(
        AHB_IF_0_AHB_BUSY), .B(N_349), .C(N_272), .D(N_357), .Y(
        un1_addr_temp_8_sqmuxa_2_i_i_i_1));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[1]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[1] ), .Y(
        \data_lm[1] ));
    SLE start_envm_reg2 (.D(start_envm_reg1_net_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        start_envm_reg2_net_1));
    CFG4 #( .INIT(16'hCAC0) )  \current_state_ns_0_0[12]  (.A(
        \current_state[11]_net_1 ), .B(\current_state[12]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_514), .Y(\current_state_ns[12] ));
    CFG4 #( .INIT(16'hA0CC) )  \addr_temp_lm_0[17]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\addr_temp_s[17] ), .C(
        \data_13[6] ), .D(N_822), .Y(\addr_temp_lm[17] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[8]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[8]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[7]_net_1 ), .S(\data_s[8] ), .Y(), .FCO(
        \data_cry[8]_net_1 ));
    SLE start_esram_reg (.D(start_esram_c), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        start_esram_reg_net_1));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[18]  (.A(N_822), .B(
        \addr_temp_s[18] ), .Y(\addr_temp_lm[18] ));
    SLE \ram_wdata[14]  (.D(AHB_IF_0_DATAOUT[14]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[14]));
    CFG4 #( .INIT(16'h1000) )  WRITE_RNO_2 (.A(
        \current_state[4]_net_1 ), .B(N_349), .C(N_516), .D(N_333), .Y(
        N_410));
    CFG4 #( .INIT(16'h0100) )  un1_current_state_20_i_0_0_a2_0_2 (.A(
        \current_state[8]_net_1 ), .B(\current_state[16]_net_1 ), .C(
        \data_13[31] ), .D(un1_current_state_20_i_0_0_a2_0_0_net_1), 
        .Y(un1_current_state_20_i_0_0_a2_0_2_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE \data[31]  (.D(\data_lm[31] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[31]));
    SLE \ram_wdata[28]  (.D(AHB_IF_0_DATAOUT[28]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[28]));
    SLE \data[8]  (.D(\data_lm[8] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[8]));
    SLE \data[26]  (.D(\data_lm[26] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[26]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[26]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[26]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[25]_net_1 ), .S(\data_s[26] ), .Y(), .FCO(
        \data_cry[26]_net_1 ));
    CFG4 #( .INIT(16'h0ACC) )  \addr_temp_lm_0[7]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\addr_temp_s[7] ), .C(
        \addr_temp_lm_0_1[7]_net_1 ), .D(N_822), .Y(\addr_temp_lm[7] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[29]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[29]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[28]_net_1 ), .S(\addr_temp_s[29] ), .Y(), .FCO(
        \addr_temp_cry[29]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \data_lm_0[12]  (.A(\data_s[12] ), .B(
        \data_13[6] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[12] ));
    CFG4 #( .INIT(16'h0008) )  WRITE_RNO_1 (.A(
        un1_current_state_16_0_0_i_0_0_a2_1_0), .B(N_516), .C(
        \current_state[2]_net_1 ), .D(\current_state[4]_net_1 ), .Y(
        un1_current_state_16_0_0_i_0_0_a2_1_2));
    CFG4 #( .INIT(16'h2333) )  WRITE_RNO_3 (.A(
        \current_state[3]_net_1 ), .B(N_531), .C(N_532), .D(N_407_2), 
        .Y(N_393_i_1));
    SLE \ram_wdata[12]  (.D(AHB_IF_0_DATAOUT[12]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[12]));
    SLE \ram_waddr[1]  (.D(N_372_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(ram_waddre), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_ram_waddr[1]));
    CFG4 #( .INIT(16'hF444) )  \current_state_RNIP0FE3[4]  (.A(N_349), 
        .B(N_370_i_i_0_a2_1_3), .C(\current_state[4]_net_1 ), .D(
        AHB_IF_0_DATAOUT[0]), .Y(N_370_i_i_0_0));
    SLE \current_state[13]  (.D(N_340_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[20]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[20]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[19]_net_1 ), .S(\data_s[20] ), .Y(), .FCO(
        \data_cry[20]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[20]  (.A(\data_s[20] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[20] ));
    CFG4 #( .INIT(16'h5FCC) )  \addr_temp_lm_0[29]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\addr_temp_s[29] ), .C(
        \data_13[6] ), .D(N_822), .Y(\addr_temp_lm[29] ));
    SLE \ram_wdata[26]  (.D(AHB_IF_0_DATAOUT[26]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[26]));
    CFG4 #( .INIT(16'h22F0) )  \data_lm_0[27]  (.A(
        \current_state[7]_net_1 ), .B(AHB_IF_0_AHB_BUSY), .C(
        \data_s[27] ), .D(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[27] ));
    CFG3 #( .INIT(8'h06) )  \data_cnt_RNO[1]  (.A(\data_cnt[1]_net_1 ), 
        .B(\data_cnt[0]_net_1 ), .C(N_314), .Y(N_320_i_0));
    CFG4 #( .INIT(16'h0400) )  \current_state_ns_i_i_0_a2[1]  (.A(
        start_envm_reg1_net_1), .B(start_envm_reg2_net_1), .C(
        esram_select_net_1), .D(\current_state[0]_net_1 ), .Y(N_461));
    CFG3 #( .INIT(8'hCE) )  \current_state_ns_0_0[16]  (.A(
        \current_state[15]_net_1 ), .B(N_439), .C(N_341), .Y(
        \current_state_ns[16] ));
    CFG2 #( .INIT(4'hE) )  \current_state_RNIHICS[7]  (.A(N_355), .B(
        \current_state[7]_net_1 ), .Y(N_314));
    CFG3 #( .INIT(8'hCA) )  \data_lm_0[5]  (.A(\data_s[5] ), .B(
        \data_13[6] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[5] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[4]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[3]_net_1 ), .S(\addr_temp_s[4] ), .Y(), .FCO(
        \addr_temp_cry[4]_net_1 ));
    SLE \addr_temp[2]  (.D(\addr_temp_lm[2] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[2]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[4]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[4]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[3]_net_1 ), .S(\data_s[4] ), .Y(), .FCO(
        \data_cry[4]_net_1 ));
    SLE \data[7]  (.D(\data_lm[7] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[7]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[25]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[25]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[24]_net_1 ), .S(\addr_temp_s[25] ), .Y(), .FCO(
        \addr_temp_cry[25]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3 (.A(
        eSRAM_eNVM_RW_0_ram_waddr[3]), .B(eSRAM_eNVM_RW_0_ram_waddr[1])
        , .C(\current_state[14]_net_1 ), .D(
        eSRAM_eNVM_RW_0_ram_waddr[4]), .Y(
        un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3_net_1));
    CFG4 #( .INIT(16'h55C3) )  \ram_waddr_RNO[3]  (.A(
        \current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ram_waddr[3]), 
        .C(N_352), .D(N_384), .Y(N_374_i_0));
    CFG4 #( .INIT(16'h7F70) )  \current_state_ns_0_0_o2_RNI27Q61[3]  (
        .A(AHB_IF_0_DATAOUT[2]), .B(AHB_IF_0_DATAOUT[1]), .C(
        \current_state[4]_net_1 ), .D(N_333), .Y(N_335));
    SLE \data[14]  (.D(\data_lm[14] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[14]));
    SLE \data[0]  (.D(\data_lm[0] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[0]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[9]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[8]_net_1 ), .S(\addr_temp_s[9] ), .Y(), .FCO(
        \addr_temp_cry[9]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[22]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[22] ), .Y(
        \data_lm[22] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[5]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[5]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[4]_net_1 ), .S(\data_s[5] ), .Y(), .FCO(
        \data_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0031) )  un1_READ_1_sqmuxa_2_i_0_a3_2 (.A(
        \current_state[8]_net_1 ), .B(\current_state[12]_net_1 ), .C(
        AHB_IF_0_DATAOUT[0]), .D(\current_state[9]_net_1 ), .Y(
        un1_READ_1_sqmuxa_2_i_0_a3_2_net_1));
    CFG4 #( .INIT(16'h0004) )  ram_wdata_0_sqmuxa_i_a6_1_4 (.A(
        \current_state[9]_net_1 ), .B(
        ram_wdata_0_sqmuxa_i_a6_1_3_net_1), .C(
        \current_state[15]_net_1 ), .D(\current_state[11]_net_1 ), .Y(
        ram_wdata_0_sqmuxa_i_a6_1_4_net_1));
    SLE \ram_waddr[3]  (.D(N_374_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(ram_waddre), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_ram_waddr[3]));
    CFG4 #( .INIT(16'hFF0E) )  \current_state_RNI6JBF1[6]  (.A(
        \current_state[6]_net_1 ), .B(\current_state[11]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_314), .Y(
        \current_state_RNI6JBF1[6]_net_1 ));
    SLE \data_cnt[3]  (.D(N_322_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        \current_state_RNI6JBF1[6]_net_1 ), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h8F80) )  \addr_temp_lm_0[11]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(\current_state[9]_net_1 ), 
        .C(N_822), .D(\addr_temp_s[11] ), .Y(\addr_temp_lm[11] ));
    CFG3 #( .INIT(8'h08) )  un1_current_state_19_i_0_0_a2_2_0 (.A(
        N_516), .B(N_335), .C(N_349), .Y(N_407_2));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[31]  (.A(\data_s[31]_net_1 ), 
        .B(\current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[31] ));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[26]  (.A(N_822), .B(
        \addr_temp_s[26] ), .Y(\addr_temp_lm[26] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[19]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[19]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[18]_net_1 ), .S(\addr_temp_s[19] ), .Y(), .FCO(
        \addr_temp_cry[19]_net_1 ));
    CFG2 #( .INIT(4'hB) )  READ32_i_0_o2_0_o6_i_o2 (.A(
        AHB_IF_0_AHB_BUSY), .B(AHB_IF_0_VALID), .Y(N_341));
    SLE \ram_wdata[13]  (.D(AHB_IF_0_DATAOUT[13]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[13]));
    CFG3 #( .INIT(8'hFE) )  \current_state_RNIKLCS[6]  (.A(
        \current_state[11]_net_1 ), .B(\current_state[5]_net_1 ), .C(
        \current_state[6]_net_1 ), .Y(N_349));
    SLE \ram_wdata[3]  (.D(AHB_IF_0_DATAOUT[3]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[3]));
    SLE \data_cnt[0]  (.D(N_453), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(\current_state_RNI6JBF1[6]_net_1 ), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \data_cnt[0]_net_1 ));
    SLE \current_state[12]  (.D(\current_state_ns[12] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[6]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[5]_net_1 ), .S(\addr_temp_s[6] ), .Y(), .FCO(
        \addr_temp_cry[6]_net_1 ));
    CFG4 #( .INIT(16'hFCFE) )  \addr_temp_cnst_i_a2_i_0_o2[5]  (.A(
        \addr_temp_cnst_i_a2_0_i_a2_0_0[8]_net_1 ), .B(N_337), .C(
        \current_state[1]_net_1 ), .D(AHB_IF_0_AHB_BUSY), .Y(N_379));
    SLE \data[15]  (.D(\data_lm[15] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[15]));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[13]  (.A(N_822), .B(
        \addr_temp_s[13] ), .Y(\addr_temp_lm[13] ));
    CFG3 #( .INIT(8'hAC) )  \data_lm_0[11]  (.A(\data_13[7] ), .B(
        \data_s[11] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[11] ));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[20]  (.A(N_822), .B(
        \addr_temp_s[20] ), .Y(\addr_temp_lm[20] ));
    CFG4 #( .INIT(16'h000D) )  \addr_temp_lm_0_1[7]  (.A(
        \current_state[5]_net_1 ), .B(AHB_IF_0_AHB_BUSY), .C(
        \current_state[9]_net_1 ), .D(N_337), .Y(
        \addr_temp_lm_0_1[7]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \current_state_RNIHJVS3[2]  (.A(
        un1_READ6_3_0_0_0_2), .B(N_337), .C(N_498), .D(N_499), .Y(
        \current_state_RNIHJVS3[2]_net_1 ));
    CFG3 #( .INIT(8'hF7) )  \current_state_ns_i_i_0_o2_0[4]  (.A(
        AHB_IF_0_DATAOUT[2]), .B(AHB_IF_0_DATAOUT[1]), .C(
        AHB_IF_0_DATAOUT[0]), .Y(N_360));
    SLE \ram_wdata[25]  (.D(AHB_IF_0_DATAOUT[25]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[25]));
    SLE \data[29]  (.D(\data_lm[29] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[29]));
    ARI1 #( .INIT(20'h4AA00) )  data_s_71 (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[0]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(data_s_71_FCO));
    CFG3 #( .INIT(8'hCA) )  \data_lm_0[6]  (.A(\data_s[6] ), .B(
        \data_13[6] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[6] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[7]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[7]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[6]_net_1 ), .S(\data_s[7] ), .Y(), .FCO(
        \data_cry[7]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \current_state_ns_0_0_o2[3]  (.A(
        AHB_IF_0_DATAOUT[0]), .B(\current_state[2]_net_1 ), .Y(N_333));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[25]  (.A(N_822), .B(
        \addr_temp_s[25] ), .Y(\addr_temp_lm[25] ));
    CFG3 #( .INIT(8'hDC) )  \data_cnst_o5_0[7]  (.A(AHB_IF_0_AHB_BUSY), 
        .B(\data_13[6] ), .C(\current_state[7]_net_1 ), .Y(
        \data_13[7] ));
    CFG3 #( .INIT(8'h01) )  un1_current_state_20_i_0_0_a2_3 (.A(
        AHB_IF_0_VALID), .B(\current_state[2]_net_1 ), .C(
        \current_state[4]_net_1 ), .Y(N_511));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[11]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[11]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[10]_net_1 ), .S(\data_s[11] ), .Y(), .FCO(
        \data_cry[11]_net_1 ));
    SLE \data[16]  (.D(\data_lm[16] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[16]));
    CFG2 #( .INIT(4'h1) )  un1_current_state_20_i_0_0_a2_0_0 (.A(
        \current_state[14]_net_1 ), .B(\current_state[3]_net_1 ), .Y(
        un1_current_state_20_i_0_0_a2_0_0_net_1));
    SLE \ram_wdata[20]  (.D(AHB_IF_0_DATAOUT[20]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[20]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[15]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[15]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[14]_net_1 ), .S(\addr_temp_s[15] ), .Y(), .FCO(
        \addr_temp_cry[15]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[31]  (.A(N_822), .B(
        \addr_temp_s[31]_net_1 ), .Y(\addr_temp_lm[31] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[8]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[7]_net_1 ), .S(\addr_temp_s[8] ), .Y(), .FCO(
        \addr_temp_cry[8]_net_1 ));
    SLE \ram_wdata[29]  (.D(AHB_IF_0_DATAOUT[29]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[29]));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[16]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[16] ), .Y(
        \data_lm[16] ));
    CFG4 #( .INIT(16'hFFFE) )  
        un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_RNIRRA81 (.A(
        \current_state[9]_net_1 ), .B(N_355), .C(N_292), .D(N_103), .Y(
        ram_waddre));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[22]  (.A(N_822), .B(
        \addr_temp_s[22] ), .Y(\addr_temp_lm[22] ));
    CFG4 #( .INIT(16'h0B00) )  \current_state_ns_0_0_a2_0[0]  (.A(
        start_envm_reg1_net_1), .B(start_envm_reg2_net_1), .C(
        esram_select_net_1), .D(\current_state[0]_net_1 ), .Y(N_465));
    SLE start_envm_reg1 (.D(state[0]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        start_envm_reg1_net_1));
    CFG4 #( .INIT(16'hF0F1) )  \current_state_RNIERJP1[6]  (.A(
        \current_state[6]_net_1 ), .B(\current_state[11]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_340), .Y(N_822));
    CFG2 #( .INIT(4'hB) )  ram_waddr_n3_0_o2 (.A(N_343), .B(
        eSRAM_eNVM_RW_0_ram_waddr[2]), .Y(N_352));
    CFG4 #( .INIT(16'h000E) )  un1_READ_1_sqmuxa_2_i_0_0 (.A(
        AHB_IF_0_AHB_BUSY), .B(un1_READ_1_sqmuxa_2_i_0_a3_2_2_net_1), 
        .C(\current_state[1]_net_1 ), .D(\current_state[14]_net_1 ), 
        .Y(un1_READ_1_sqmuxa_2_i_0_0_net_1));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[21]  (.A(\data_s[21] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[21] ));
    SLE \addr_temp[14]  (.D(\addr_temp_lm[14] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[14]));
    CFG4 #( .INIT(16'h0010) )  \current_state_RNI2FBF1[16]  (.A(
        \current_state[0]_net_1 ), .B(\current_state[16]_net_1 ), .C(
        un1_current_state_16_0_0_i_0_0_a2_2_0), .D(\data_13[31] ), .Y(
        N_530));
    CFG3 #( .INIT(8'h80) )  \current_state_ns_0_0_a2_0[16]  (.A(
        envm_release_reg_net_1), .B(\current_state[16]_net_1 ), .C(
        AHB_IF_0_AHB_BUSY), .Y(N_439));
    SLE \current_state[7]  (.D(\current_state_ns[7] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[13]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[13]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[12]_net_1 ), .S(\data_s[13] ), .Y(), .FCO(
        \data_cry[13]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  un1_ram_wen_0_sqmuxa_i_0_0_0 (.A(
        \current_state[9]_net_1 ), .B(N_355), .C(N_103), .Y(N_384));
    CFG4 #( .INIT(16'hF1F0) )  un1_current_state_20_i_0_0_0 (.A(
        \current_state[1]_net_1 ), .B(\current_state[14]_net_1 ), .C(
        N_448), .D(N_530), .Y(un1_current_state_20_i_0_0_0_net_1));
    SLE READ (.D(N_379_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        N_391_i_0), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(eSRAM_eNVM_RW_0_READ));
    CFG3 #( .INIT(8'hCA) )  \data_lm_0[4]  (.A(\data_s[4] ), .B(
        \data_13[6] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[4] ));
    CFG4 #( .INIT(16'h0CAE) )  \current_state_ns_0[8]  (.A(
        \current_state[7]_net_1 ), .B(\current_state[8]_net_1 ), .C(
        AHB_IF_0_DATAOUT[0]), .D(AHB_IF_0_AHB_BUSY), .Y(
        \current_state_ns[8] ));
    SLE \addr_temp[24]  (.D(\addr_temp_lm[24] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[24]));
    SLE \data[2]  (.D(\data_lm[2] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[2]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[2]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[2]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[1]_net_1 ), .S(\data_s[2] ), .Y(), .FCO(
        \data_cry[2]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \current_state_RNI6AUF[16]  (.A(
        \current_state[7]_net_1 ), .B(\data_13[31] ), .C(
        \current_state[16]_net_1 ), .Y(N_516));
    SLE ram_wen (.D(N_292), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        N_388_i_0), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(eSRAM_eNVM_RW_0_ram_wen));
    SLE \addr_temp[4]  (.D(\addr_temp_lm[4] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[4]));
    CFG4 #( .INIT(16'h0203) )  
        un1_current_state_19_i_0_0_a2_2_0_RNI1K2N5 (.A(
        \current_state[0]_net_1 ), .B(N_530), .C(N_370_i_i_0_0), .D(
        N_407_2), .Y(N_141_i_0));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[26]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[26] ), .Y(
        \data_lm[26] ));
    CFG3 #( .INIT(8'hE0) )  \current_state_RNIKLCS[2]  (.A(
        \current_state[4]_net_1 ), .B(\current_state[2]_net_1 ), .C(
        \current_state[16]_net_1 ), .Y(N_498));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[21]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[21]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[20]_net_1 ), .S(\data_s[21] ), .Y(), .FCO(
        \data_cry[21]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[23]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[23]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[22]_net_1 ), .S(\addr_temp_s[23] ), .Y(), .FCO(
        \addr_temp_cry[23]_net_1 ));
    SLE \data[27]  (.D(\data_lm[27] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[27]));
    CFG4 #( .INIT(16'hECA0) )  envm_release_reg_RNI8QJR (.A(
        envm_release_reg_net_1), .B(\current_state[2]_net_1 ), .C(
        \current_state[16]_net_1 ), .D(AHB_IF_0_DATAOUT[0]), .Y(N_337));
    CFG3 #( .INIT(8'h0E) )  \current_state_RNIEA38[15]  (.A(
        \current_state[15]_net_1 ), .B(\current_state[14]_net_1 ), .C(
        N_341), .Y(N_292));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_s[31]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[31]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[30]_net_1 ), .S(\addr_temp_s[31]_net_1 ), .Y(), 
        .FCO());
    CFG2 #( .INIT(4'h4) )  \addr_temp_cnst_i_a2_0_i_a2_0_0[8]  (.A(
        AHB_IF_0_DATAOUT[0]), .B(\current_state[8]_net_1 ), .Y(
        \addr_temp_cnst_i_a2_0_i_a2_0_0[8]_net_1 ));
    SLE \ram_wdata[27]  (.D(AHB_IF_0_DATAOUT[27]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[27]));
    CFG3 #( .INIT(8'h15) )  WRITE_RNO_7 (.A(\current_state[2]_net_1 ), 
        .B(AHB_IF_0_DATAOUT[2]), .C(AHB_IF_0_DATAOUT[1]), .Y(
        un1_current_state_16_0_0_i_0_0_a2_0_0));
    SLE \data[28]  (.D(\data_lm[28] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[28]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[3]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[3]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[2]_net_1 ), .S(\data_s[3] ), .Y(), .FCO(
        \data_cry[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  esram_select (.A(start_esram_reg1_net_1), 
        .B(start_esram_reg2_net_1), .Y(esram_select_net_1));
    CFG4 #( .INIT(16'h2C2E) )  \current_state_RNO[11]  (.A(
        \current_state[11]_net_1 ), .B(\data_13[31] ), .C(
        AHB_IF_0_AHB_BUSY), .D(N_514), .Y(N_337_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[12]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[12]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[11]_net_1 ), .S(\data_s[12] ), .Y(), .FCO(
        \data_cry[12]_net_1 ));
    CFG2 #( .INIT(4'hB) )  ram_waddr_n4_0_o2 (.A(N_352), .B(
        eSRAM_eNVM_RW_0_ram_waddr[3]), .Y(N_362));
    SLE envm_release_reg (.D(\current_state[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un40_0_0_0_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        envm_release_reg_net_1));
    CFG4 #( .INIT(16'h03A3) )  \addr_temp_lm_0[2]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(eSRAM_eNVM_RW_0_ADDR[2]), 
        .C(N_822), .D(\addr_temp_lm_0_1_0[2]_net_1 ), .Y(
        \addr_temp_lm[2] ));
    CFG4 #( .INIT(16'hFC55) )  \data_lm_0[0]  (.A(
        eSRAM_eNVM_RW_0_DATAOUT[0]), .B(\data_lm_0_1_0[0]_net_1 ), .C(
        \data_13[6] ), .D(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[0] ));
    CFG2 #( .INIT(4'h1) )  un1_current_state_13_i_0_0_a2_0 (.A(
        \current_state[16]_net_1 ), .B(\current_state[13]_net_1 ), .Y(
        un1_current_state_13_i_0_0_a2_0_net_1));
    SLE \data[19]  (.D(\data_lm[19] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[19]));
    CFG4 #( .INIT(16'h0001) )  ram_wdata_0_sqmuxa_i_a6_1_3 (.A(
        \current_state[1]_net_1 ), .B(\current_state[7]_net_1 ), .C(
        \current_state[3]_net_1 ), .D(\current_state[5]_net_1 ), .Y(
        ram_wdata_0_sqmuxa_i_a6_1_3_net_1));
    SLE \ram_waddr[0]  (.D(N_9_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(ram_waddre), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_ram_waddr[0]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[23]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[23]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[22]_net_1 ), .S(\data_s[23] ), .Y(), .FCO(
        \data_cry[23]_net_1 ));
    SLE \current_state[4]  (.D(\current_state_ns_i_i_0[4]_net_1 ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[4]_net_1 ));
    SLE \data[22]  (.D(\data_lm[22] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[22]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[30]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[30]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[29]_net_1 ), .S(\addr_temp_s[30] ), .Y(), .FCO(
        \addr_temp_cry[30]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \data_lm_0[7]  (.A(\data_13[7] ), .B(
        \data_s[7] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .Y(
        \data_lm[7] ));
    SLE \addr_temp[10]  (.D(\addr_temp_lm[10] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[10]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[15]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[15]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[14]_net_1 ), .S(\data_s[15] ), .Y(), .FCO(
        \data_cry[15]_net_1 ));
    SLE \ram_waddr[2]  (.D(N_373_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(ram_waddre), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_ram_waddr[2]));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[14]  (.A(N_822), .B(
        \addr_temp_s[14] ), .Y(\addr_temp_lm[14] ));
    SLE \addr_temp[8]  (.D(\addr_temp_lm[8] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[8]));
    ARI1 #( .INIT(20'h4AA00) )  \data_s[31]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[31]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[30]_net_1 ), .S(\data_s[31]_net_1 ), .Y(), .FCO(
        ));
    CFG4 #( .INIT(16'h44AE) )  \current_state_RNO[6]  (.A(
        \current_state[5]_net_1 ), .B(\current_state[6]_net_1 ), .C(
        N_514), .D(AHB_IF_0_AHB_BUSY), .Y(N_331_i_0));
    SLE \current_state[10]  (.D(\current_state_ns[10] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\data_13[31] ));
    SLE \current_state[0]  (.D(\current_state_ns[0] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[0]_net_1 ));
    SLE \ram_wdata[18]  (.D(AHB_IF_0_DATAOUT[18]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[18]));
    SLE \addr_temp[9]  (.D(\addr_temp_lm[9] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[9]));
    SLE \ram_wdata[7]  (.D(AHB_IF_0_DATAOUT[7]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[7]));
    SLE \addr_temp[20]  (.D(\addr_temp_lm[20] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[20]));
    SLE \addr_temp[17]  (.D(\addr_temp_lm[17] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[17]));
    SLE \addr_temp[5]  (.D(\addr_temp_lm[5] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[5]));
    CFG4 #( .INIT(16'hF4F0) )  \current_state_ns_i_i_0[1]  (.A(
        \current_state[0]_net_1 ), .B(\current_state[1]_net_1 ), .C(
        N_461), .D(AHB_IF_0_AHB_BUSY), .Y(
        \current_state_ns_i_i_0[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[13]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[12]_net_1 ), .S(\addr_temp_s[13] ), .Y(), .FCO(
        \addr_temp_cry[13]_net_1 ));
    SLE \addr_temp[11]  (.D(\addr_temp_lm[11] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[11]));
    CFG4 #( .INIT(16'h5501) )  ram_wdata_0_sqmuxa_i_a6_1_4_RNI4B9G1 (
        .A(ram_wdata_0_sqmuxa_i_0_net_1), .B(
        ram_wdata_0_sqmuxa_i_a6_1_4_net_1), .C(
        ram_wdata_0_sqmuxa_i_2_tz_net_1), .D(N_340), .Y(N_149_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[28]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[28]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[27]_net_1 ), .S(\addr_temp_s[28] ), .Y(), .FCO(
        \addr_temp_cry[28]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[1]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[1]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(data_s_71_FCO), .S(\data_s[1] ), .Y(), .FCO(
        \data_cry[1]_net_1 ));
    CFG3 #( .INIT(8'h10) )  un1_current_state_20_i_0_0_a2_4 (.A(
        \current_state[13]_net_1 ), .B(\current_state[9]_net_1 ), .C(
        N_335), .Y(N_512));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[27]  (.A(N_822), .B(
        \addr_temp_s[27] ), .Y(\addr_temp_lm[27] ));
    SLE \ram_wdata[2]  (.D(AHB_IF_0_DATAOUT[2]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[2]));
    CFG3 #( .INIT(8'hF2) )  \addr_temp_cnst_i_a2_0_i_o2_1_0[8]  (.A(
        \current_state[7]_net_1 ), .B(AHB_IF_0_AHB_BUSY), .C(
        \current_state[1]_net_1 ), .Y(
        \addr_temp_cnst_i_a2_0_i_o2_1_0[8]_net_1 ));
    SLE \addr_temp[27]  (.D(\addr_temp_lm[27] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[27]));
    SLE \ram_wdata[16]  (.D(AHB_IF_0_DATAOUT[16]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[16]));
    CFG2 #( .INIT(4'hB) )  ram_wdata_0_sqmuxa_i_0 (.A(N_341), .B(
        eSRAM_eNVM_access_0_HPMS_READY), .Y(
        ram_wdata_0_sqmuxa_i_0_net_1));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[28]  (.A(N_822), .B(
        \addr_temp_s[28] ), .Y(\addr_temp_lm[28] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[22]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[22]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[21]_net_1 ), .S(\data_s[22] ), .Y(), .FCO(
        \data_cry[22]_net_1 ));
    SLE \addr_temp[21]  (.D(\addr_temp_lm[21] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[21]));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[14]  (.A(\data_s[14] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[14] ));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[5]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[4]_net_1 ), .S(\addr_temp_s[5] ), .Y(), .FCO(
        \addr_temp_cry[5]_net_1 ));
    SLE \current_state[14]  (.D(N_342_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[14]_net_1 ));
    SLE \addr_temp[19]  (.D(\addr_temp_lm[19] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[19]));
    SLE \ram_wdata[21]  (.D(AHB_IF_0_DATAOUT[21]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[21]));
    SLE \current_state[11]  (.D(N_337_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[11]_net_1 ));
    CFG4 #( .INIT(16'hCA0A) )  \addr_temp_lm_0[6]  (.A(
        \addr_temp_s[6] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_241), .Y(\addr_temp_lm[6] ));
    CFG4 #( .INIT(16'hAAAE) )  WRITE_RNO_6 (.A(N_531), .B(
        un1_current_state_16_0_0_i_0_0_a2_2_0), .C(
        \current_state[16]_net_1 ), .D(\data_13[31] ), .Y(
        un1_current_state_16_0_0_i_0_0_0));
    CFG2 #( .INIT(4'h4) )  \data_lm_0[19]  (.A(
        \current_state_RNIHJVS3[2]_net_1 ), .B(\data_s[19] ), .Y(
        \data_lm[19] ));
    CFG4 #( .INIT(16'h0001) )  envm_release_reg_RNIKPH21 (.A(
        \current_state[7]_net_1 ), .B(envm_release_reg_net_1), .C(
        \data_13[31] ), .D(\current_state[0]_net_1 ), .Y(
        N_370_i_i_0_a2_1_2));
    CFG4 #( .INIT(16'hCA0A) )  \addr_temp_lm_0[5]  (.A(
        \addr_temp_s[5] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_379), .Y(\addr_temp_lm[5] ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[25]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[25]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[24]_net_1 ), .S(\data_s[25] ), .Y(), .FCO(
        \data_cry[25]_net_1 ));
    SLE \data[17]  (.D(\data_lm[17] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[17]));
    SLE \addr_temp[29]  (.D(\addr_temp_lm[29] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[29]));
    CFG2 #( .INIT(4'h4) )  \data_cnst_o5_0_a2_0_a2[8]  (.A(N_360), .B(
        \current_state[4]_net_1 ), .Y(\data_13[6] ));
    SLE \current_state[8]  (.D(\current_state_ns[8] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[8]_net_1 ));
    SLE \current_state[1]  (.D(\current_state_ns_i_i_0[1]_net_1 ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[1]_net_1 ));
    SLE \current_state[15]  (.D(\current_state_ns[15] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[15]_net_1 ));
    CFG4 #( .INIT(16'h5595) )  data_cnt_n4_i_x2 (.A(
        \data_cnt[4]_net_1 ), .B(\data_cnt[3]_net_1 ), .C(
        \data_cnt[2]_net_1 ), .D(N_339), .Y(N_347_i));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[21]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[21]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[20]_net_1 ), .S(\addr_temp_s[21] ), .Y(), .FCO(
        \addr_temp_cry[21]_net_1 ));
    SLE WRITE (.D(N_793_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        N_393_i_0), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(eSRAM_eNVM_RW_0_WRITE));
    CFG2 #( .INIT(4'h1) )  \data_cnt_RNO[4]  (.A(N_314), .B(N_347_i), 
        .Y(N_323_i_0));
    SLE \data[18]  (.D(\data_lm[18] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[18]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[14]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[14]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[13]_net_1 ), .S(\data_s[14] ), .Y(), .FCO(
        \data_cry[14]_net_1 ));
    SLE \data[20]  (.D(\data_lm[20] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[20]));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[22]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[22]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[21]_net_1 ), .S(\addr_temp_s[22] ), .Y(), .FCO(
        \addr_temp_cry[22]_net_1 ));
    SLE \current_state[3]  (.D(\current_state_ns[3] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[3]_net_1 ));
    CFG4 #( .INIT(16'h440C) )  
        \addr_temp_cnst_0_a2_i_0_o2_1_RNI26573[19]  (.A(N_341), .B(
        eSRAM_eNVM_access_0_HPMS_READY), .C(
        un1_addr_temp_8_sqmuxa_2_i_i_i_1), .D(N_340), .Y(N_40));
    CFG4 #( .INIT(16'h5554) )  \current_state_RNO[13]  (.A(
        \current_state_ns_i_0_0_0[13]_net_1 ), .B(N_341), .C(
        \current_state[12]_net_1 ), .D(\current_state[9]_net_1 ), .Y(
        N_340_i_0));
    SLE \current_state[9]  (.D(\current_state_ns[9] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \current_state[9]_net_1 ));
    SLE \data[23]  (.D(\data_lm[23] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[23]));
    CFG3 #( .INIT(8'hC5) )  \current_state_ns_0_0[3]  (.A(N_333), .B(
        \current_state[3]_net_1 ), .C(AHB_IF_0_AHB_BUSY), .Y(
        \current_state_ns[3] ));
    CFG4 #( .INIT(16'hCCEC) )  WRITE_RNO_4 (.A(N_516), .B(
        un1_current_state_16_0_0_i_0_0_0), .C(
        un1_current_state_16_0_0_i_0_0_a2_0_0), .D(N_349), .Y(
        un1_current_state_16_0_0_i_0_0_1));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[18]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[18]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[17]_net_1 ), .S(\addr_temp_s[18] ), .Y(), .FCO(
        \addr_temp_cry[18]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[24]  (.A(\data_s[24] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[24] ));
    CFG3 #( .INIT(8'h04) )  \current_state_RNIK3PT1[2]  (.A(
        \current_state[4]_net_1 ), .B(N_370_i_i_0_a2_1_2), .C(
        \current_state[2]_net_1 ), .Y(N_370_i_i_0_a2_1_3));
    CFG4 #( .INIT(16'h0054) )  WRITE_RNO_0 (.A(N_448), .B(
        \current_state[8]_net_1 ), .C(N_393_i_1), .D(N_409), .Y(
        N_393_i_0));
    CFG4 #( .INIT(16'h0F0D) )  ram_wen_RNO (.A(
        un1_current_state_13_i_0_0_a2_0_net_1), .B(
        \current_state[0]_net_1 ), .C(N_103), .D(N_292), .Y(N_388_i_0));
    CFG3 #( .INIT(8'hE2) )  \data_lm_0[29]  (.A(\data_s[29] ), .B(
        \current_state_RNIHJVS3[2]_net_1 ), .C(\data_13[31] ), .Y(
        \data_lm[29] ));
    CFG4 #( .INIT(16'h3AFA) )  \addr_temp_lm_0[19]  (.A(
        \addr_temp_s[19] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_272), .Y(\addr_temp_lm[19] ));
    CFG3 #( .INIT(8'hAE) )  \addr_temp_cnst_i_a2_i_a6_0_o2[6]  (.A(
        N_337), .B(\current_state[7]_net_1 ), .C(AHB_IF_0_AHB_BUSY), 
        .Y(N_241));
    CFG4 #( .INIT(16'hFACA) )  \data_lm_0[9]  (.A(\data_s[9] ), .B(
        \data_13[31] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .D(
        \data_13[6] ), .Y(\data_lm[9] ));
    SLE \addr_temp[12]  (.D(\addr_temp_lm[12] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[12]));
    SLE \ram_wdata[24]  (.D(AHB_IF_0_DATAOUT[24]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[24]));
    CFG4 #( .INIT(16'hEAC0) )  \current_state_ns_0_0[10]  (.A(
        AHB_IF_0_AHB_BUSY), .B(esram_select_net_1), .C(
        \current_state[0]_net_1 ), .D(\data_13[31] ), .Y(
        \current_state_ns[10] ));
    CFG4 #( .INIT(16'hFACA) )  \data_lm_0[8]  (.A(\data_s[8] ), .B(
        \data_13[31] ), .C(\current_state_RNIHJVS3[2]_net_1 ), .D(
        \data_13[6] ), .Y(\data_lm[8] ));
    SLE \data[12]  (.D(\data_lm[12] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[12]));
    SLE \addr_temp[18]  (.D(\addr_temp_lm[18] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[18]));
    CFG4 #( .INIT(16'h0007) )  READ_RNO (.A(
        un1_READ_1_sqmuxa_2_i_0_a3_2_net_1), .B(
        un1_READ_1_sqmuxa_2_i_0_a3_1_net_1), .C(N_103), .D(
        un1_READ_1_sqmuxa_2_i_0_0_net_1), .Y(N_379_i_0));
    SLE \ram_wdata[15]  (.D(AHB_IF_0_DATAOUT[15]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[15]));
    SLE \ram_wdata[1]  (.D(AHB_IF_0_DATAOUT[1]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[1]));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[19]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[19]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[18]_net_1 ), .S(\data_s[19] ), .Y(), .FCO(
        \data_cry[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[18]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[18]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[17]_net_1 ), .S(\data_s[18] ), .Y(), .FCO(
        \data_cry[18]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \data_cry[30]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_DATAOUT[30]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\data_cry[29]_net_1 ), .S(\data_s[30] ), .Y(), .FCO(
        \data_cry[30]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \current_state_RNI4SUQ[4]  (.A(
        AHB_IF_0_DATAOUT[1]), .B(\current_state[4]_net_1 ), .C(
        AHB_IF_0_DATAOUT[2]), .Y(N_499));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[21]  (.A(N_822), .B(
        \addr_temp_s[21] ), .Y(\addr_temp_lm[21] ));
    SLE \addr_temp[22]  (.D(\addr_temp_lm[22] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[22]));
    SLE \ram_wdata[22]  (.D(AHB_IF_0_DATAOUT[22]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[22]));
    SLE \ram_wdata[10]  (.D(AHB_IF_0_DATAOUT[10]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[10]));
    CFG4 #( .INIT(16'hCA0A) )  \addr_temp_lm_0[8]  (.A(
        \addr_temp_s[8] ), .B(eSRAM_eNVM_access_0_HPMS_READY), .C(
        N_822), .D(N_357), .Y(\addr_temp_lm[8] ));
    SLE \data[21]  (.D(\data_lm[21] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[21]));
    SLE \addr_temp[28]  (.D(\addr_temp_lm[28] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[28]));
    CFG4 #( .INIT(16'hF0F8) )  un40_0_0_0 (.A(
        \current_state[16]_net_1 ), .B(envm_release_reg_net_1), .C(
        \current_state[9]_net_1 ), .D(AHB_IF_0_AHB_BUSY), .Y(
        un40_0_0_0_net_1));
    CFG4 #( .INIT(16'h00A6) )  \data_cnt_RNO[3]  (.A(
        \data_cnt[3]_net_1 ), .B(\data_cnt[2]_net_1 ), .C(N_339), .D(
        N_314), .Y(N_322_i_0));
    CFG2 #( .INIT(4'h4) )  \addr_temp_lm_0[23]  (.A(N_822), .B(
        \addr_temp_s[23] ), .Y(\addr_temp_lm[23] ));
    SLE \addr_temp[15]  (.D(\addr_temp_lm[15] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_40), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ADDR[15]));
    CFG4 #( .INIT(16'h0001) )  ram_wdata_0_sqmuxa_i_a6_0_4_2 (.A(
        \current_state[14]_net_1 ), .B(\current_state[7]_net_1 ), .C(
        \current_state[15]_net_1 ), .D(\current_state[5]_net_1 ), .Y(
        ram_wdata_0_sqmuxa_i_a6_0_4_2_net_1));
    SLE \ram_wdata[19]  (.D(AHB_IF_0_DATAOUT[19]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[19]));
    SLE \ram_wdata[0]  (.D(AHB_IF_0_DATAOUT[0]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[0]));
    SLE \ram_wdata[30]  (.D(AHB_IF_0_DATAOUT[30]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_149_i_0), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(eSRAM_eNVM_RW_0_ram_wdata[30]));
    CFG3 #( .INIT(8'hF8) )  \current_state_ns_0[15]  (.A(
        \current_state[15]_net_1 ), .B(N_341), .C(N_103), .Y(
        \current_state_ns[15] ));
    CFG4 #( .INIT(16'hFFCE) )  
        un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3_RNIPQK61 (.A(
        \current_state[14]_net_1 ), .B(\current_state[13]_net_1 ), .C(
        un1_READ_1_sqmuxa_2_i_0_a3_0_0_a2_3_net_1), .D(
        un1_addr_temp_8_sqmuxa_2_i_i_o2_3_0_c), .Y(N_340));
    ARI1 #( .INIT(20'h4AA00) )  \addr_temp_cry[11]  (.A(VCC_net_1), .B(
        eSRAM_eNVM_RW_0_ADDR[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        \addr_temp_cry[10]_net_1 ), .S(\addr_temp_s[11] ), .Y(), .FCO(
        \addr_temp_cry[11]_net_1 ));
    SLE \data[3]  (.D(\data_lm[3] ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_141_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        eSRAM_eNVM_RW_0_DATAOUT[3]));
    
endmodule


module 
        AHB_IF_0s_1s_2s_3s_4294967292s_4294967293s_4294967294s_0s_1_layer0(
        
       eSRAM_eNVM_RW_0_DATAOUT,
       AHB_IF_0_DATAOUT,
       AHB_IF_0_BIF_1_HRDATA,
       AHB_IF_0_BIF_1_HWDATA,
       AHB_IF_0_BIF_1_HADDR,
       AHB_IF_0_BIF_1_HTRANS,
       eSRAM_eNVM_RW_0_ADDR,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       eSRAM_eNVM_access_0_HPMS_READY,
       AHB_IF_0_VALID,
       AHB_IF_0_AHB_BUSY,
       AHB_IF_0_BIF_1_HWRITE,
       HREADY_M_0_iv_i_0,
       eSRAM_eNVM_RW_0_WRITE,
       eSRAM_eNVM_RW_0_READ,
       N_546,
       defSlaveSMCurrentState,
       N_53,
       defSlaveSMNextState
    );
input  [31:0] eSRAM_eNVM_RW_0_DATAOUT;
output [31:0] AHB_IF_0_DATAOUT;
input  [31:0] AHB_IF_0_BIF_1_HRDATA;
output [31:0] AHB_IF_0_BIF_1_HWDATA;
output [31:2] AHB_IF_0_BIF_1_HADDR;
output [1:1] AHB_IF_0_BIF_1_HTRANS;
input  [31:2] eSRAM_eNVM_RW_0_ADDR;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
input  eSRAM_eNVM_access_0_HPMS_READY;
output AHB_IF_0_VALID;
output AHB_IF_0_AHB_BUSY;
output AHB_IF_0_BIF_1_HWRITE;
input  HREADY_M_0_iv_i_0;
input  eSRAM_eNVM_RW_0_WRITE;
input  eSRAM_eNVM_RW_0_READ;
input  N_546;
input  defSlaveSMCurrentState;
input  N_53;
input  defSlaveSMNextState;

    wire \HWDATA_int[20]_net_1 , VCC_net_1, N_47_i_0, GND_net_1, 
        \HWDATA_int[21]_net_1 , \HWDATA_int[22]_net_1 , 
        \HWDATA_int[23]_net_1 , \HWDATA_int[24]_net_1 , 
        \HWDATA_int[25]_net_1 , \HWDATA_int[26]_net_1 , 
        \HWDATA_int[27]_net_1 , \HWDATA_int[28]_net_1 , 
        \HWDATA_int[29]_net_1 , \HWDATA_int[30]_net_1 , 
        \HWDATA_int[31]_net_1 , \HWDATA_int[5]_net_1 , 
        \HWDATA_int[6]_net_1 , \HWDATA_int[7]_net_1 , 
        \HWDATA_int[8]_net_1 , \HWDATA_int[9]_net_1 , 
        \HWDATA_int[10]_net_1 , \HWDATA_int[11]_net_1 , 
        \HWDATA_int[12]_net_1 , \HWDATA_int[13]_net_1 , 
        \HWDATA_int[14]_net_1 , \HWDATA_int[15]_net_1 , 
        \HWDATA_int[16]_net_1 , \HWDATA_int[17]_net_1 , 
        \HWDATA_int[18]_net_1 , \HWDATA_int[19]_net_1 , 
        DATAOUT_1_sqmuxa, \HWDATA_int[0]_net_1 , \HWDATA_int[1]_net_1 , 
        \HWDATA_int[2]_net_1 , \HWDATA_int[3]_net_1 , 
        \HWDATA_int[4]_net_1 , HWDATA_1_sqmuxa, \HADDR_6[26]_net_1 , 
        N_101_i_0, \HADDR_6[27]_net_1 , \HADDR_6[28]_net_1 , 
        \HADDR_6[29]_net_1 , \HADDR_6[30]_net_1 , \HADDR_6[31]_net_1 , 
        \HADDR_6[11]_net_1 , \HADDR_6[12]_net_1 , \HADDR_6[13]_net_1 , 
        \HADDR_6[14]_net_1 , \HADDR_6[15]_net_1 , \HADDR_6[16]_net_1 , 
        \HADDR_6[17]_net_1 , \HADDR_6[18]_net_1 , \HADDR_6[19]_net_1 , 
        \HADDR_6[20]_net_1 , \HADDR_6[21]_net_1 , \HADDR_6[22]_net_1 , 
        \HADDR_6[23]_net_1 , \HADDR_6[24]_net_1 , \HADDR_6[25]_net_1 , 
        \HADDR_6[2]_net_1 , \HADDR_6[3]_net_1 , \HADDR_6[4]_net_1 , 
        \HADDR_6[5]_net_1 , \HADDR_6[6]_net_1 , \HADDR_6[7]_net_1 , 
        \HADDR_6[8]_net_1 , \HADDR_6[9]_net_1 , \HADDR_6[10]_net_1 , 
        un18_N_5_mux_i_0, N_21, N_106_i_0, N_46, un1_N_5_mux_0_i_0, 
        \ahb_fsm_current_state[1]_net_1 , un1_N_5_mux_i_0, 
        \ahb_fsm_current_state[0]_net_1 , 
        \ahb_fsm_current_state_ns[0] , N_94_i_0, 
        \ahb_fsm_current_state[2]_net_1 , 
        \ahb_fsm_current_state_ns[2] , 
        \ahb_fsm_current_state[3]_net_1 , 
        \ahb_fsm_current_state[4]_net_1 , 
        \ahb_fsm_current_state_ns[4] , 
        \ahb_fsm_current_state[5]_net_1 , 
        \ahb_fsm_current_state_ns[5] , 
        \ahb_fsm_current_state[6]_net_1 , N_115, N_52, N_84, 
        un1_m2_0_a2_0_0, N_63, N_22, un1_HADDR_0_sqmuxa_i_0_a2_c;
    
    SLE \HADDR[9]  (.D(\HADDR_6[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[9]));
    SLE \HADDR[19]  (.D(\HADDR_6[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[19]));
    SLE \DATAOUT[2]  (.D(AHB_IF_0_BIF_1_HRDATA[2]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[2]));
    SLE \HADDR[8]  (.D(\HADDR_6[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[8]));
    SLE \HWDATA_int[0]  (.D(eSRAM_eNVM_RW_0_DATAOUT[0]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[0]_net_1 ));
    SLE \HWDATA_int[29]  (.D(eSRAM_eNVM_RW_0_DATAOUT[29]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[29]_net_1 ));
    SLE \HWDATA[5]  (.D(\HWDATA_int[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[5]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[10]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[10])
        , .Y(\HADDR_6[10]_net_1 ));
    SLE \ahb_fsm_current_state[3]  (.D(
        \ahb_fsm_current_state[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HREADY_M_0_iv_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[3]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[3]), 
        .Y(\HADDR_6[3]_net_1 ));
    SLE \DATAOUT[1]  (.D(AHB_IF_0_BIF_1_HRDATA[1]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[1]));
    SLE \DATAOUT[21]  (.D(AHB_IF_0_BIF_1_HRDATA[21]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[21]));
    SLE \DATAOUT[22]  (.D(AHB_IF_0_BIF_1_HRDATA[22]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[22]));
    CFG4 #( .INIT(16'h0203) )  un1_HADDR_0_sqmuxa_i_0_o2_s_0_RNIJLTK1 
        (.A(\ahb_fsm_current_state[0]_net_1 ), .B(N_52), .C(
        un1_HADDR_0_sqmuxa_i_0_a2_c), .D(N_53), .Y(N_101_i_0));
    SLE \HWDATA_int[9]  (.D(eSRAM_eNVM_RW_0_DATAOUT[9]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[9]_net_1 ));
    SLE \ahb_fsm_current_state[5]  (.D(\ahb_fsm_current_state_ns[5] ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[5]_net_1 ));
    SLE \HADDR[6]  (.D(\HADDR_6[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[6]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[29]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[29])
        , .Y(\HADDR_6[29]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[28]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[28])
        , .Y(\HADDR_6[28]_net_1 ));
    SLE \DATAOUT[23]  (.D(AHB_IF_0_BIF_1_HRDATA[23]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[23]));
    SLE \HADDR[18]  (.D(\HADDR_6[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[18]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[5]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[5]), 
        .Y(\HADDR_6[5]_net_1 ));
    SLE \HWDATA_int[7]  (.D(eSRAM_eNVM_RW_0_DATAOUT[7]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[7]_net_1 ));
    SLE \HWDATA_int[18]  (.D(eSRAM_eNVM_RW_0_DATAOUT[18]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[18]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[27]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[27])
        , .Y(\HADDR_6[27]_net_1 ));
    SLE \HADDR[3]  (.D(\HADDR_6[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[3]));
    SLE \DATAOUT[0]  (.D(AHB_IF_0_BIF_1_HRDATA[0]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[0]));
    CFG3 #( .INIT(8'h80) )  \ahb_fsm_current_state_RNI9TCO[0]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(
        eSRAM_eNVM_access_0_HPMS_READY), .C(eSRAM_eNVM_RW_0_WRITE), .Y(
        N_47_i_0));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[15]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[15])
        , .Y(\HADDR_6[15]_net_1 ));
    SLE \DATAOUT[14]  (.D(AHB_IF_0_BIF_1_HRDATA[14]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[14]));
    SLE \DATAOUT[28]  (.D(AHB_IF_0_BIF_1_HRDATA[28]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[28]));
    SLE \HWDATA[2]  (.D(\HWDATA_int[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[2]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[30]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[30])
        , .Y(\HADDR_6[30]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[8]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[8]), 
        .Y(\HADDR_6[8]_net_1 ));
    SLE \DATAOUT[3]  (.D(AHB_IF_0_BIF_1_HRDATA[3]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[3]));
    CFG4 #( .INIT(16'h005D) )  un1_HADDR_0_sqmuxa_i_0_o2_s_0 (.A(N_22), 
        .B(N_546), .C(defSlaveSMCurrentState), .D(
        \ahb_fsm_current_state[0]_net_1 ), .Y(
        un1_HADDR_0_sqmuxa_i_0_a2_c));
    CFG2 #( .INIT(4'h8) )  \ahb_fsm_current_state_RNO[1]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_WRITE), 
        .Y(N_94_i_0));
    CFG2 #( .INIT(4'hE) )  HTRANS_2_i_o3_i_a2_0_o2 (.A(
        \ahb_fsm_current_state[2]_net_1 ), .B(
        \ahb_fsm_current_state[5]_net_1 ), .Y(N_22));
    SLE \HWDATA_int[16]  (.D(eSRAM_eNVM_RW_0_DATAOUT[16]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[16]_net_1 ));
    SLE \HADDR[29]  (.D(\HADDR_6[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[29]));
    SLE \ahb_fsm_current_state[1]  (.D(N_94_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[1]_net_1 ));
    SLE \HWDATA[3]  (.D(\HWDATA_int[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[3]));
    SLE \DATAOUT[30]  (.D(AHB_IF_0_BIF_1_HRDATA[30]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[30]));
    SLE \HWDATA_int[1]  (.D(eSRAM_eNVM_RW_0_DATAOUT[1]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \HADDR[12]  (.D(\HADDR_6[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[12]));
    CFG4 #( .INIT(16'h555D) )  \HTRANS_1_RNO[1]  (.A(un1_m2_0_a2_0_0), 
        .B(\ahb_fsm_current_state[5]_net_1 ), .C(N_53), .D(
        defSlaveSMNextState), .Y(un1_N_5_mux_0_i_0));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[14]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[14])
        , .Y(\HADDR_6[14]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  AHB_BUSY_RNO (.A(N_53), .B(
        \ahb_fsm_current_state[0]_net_1 ), .C(defSlaveSMNextState), .Y(
        N_21));
    SLE \HWDATA[17]  (.D(\HWDATA_int[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[17]));
    SLE \DATAOUT[17]  (.D(AHB_IF_0_BIF_1_HRDATA[17]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[17]));
    SLE \HADDR[28]  (.D(\HADDR_6[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[28]));
    SLE \HADDR[13]  (.D(\HADDR_6[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[13]));
    SLE \DATAOUT[26]  (.D(AHB_IF_0_BIF_1_HRDATA[26]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[26]));
    SLE AHB_BUSY (.D(N_21), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        N_106_i_0), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(AHB_IF_0_AHB_BUSY));
    SLE \ahb_fsm_current_state[4]  (.D(\ahb_fsm_current_state_ns[4] ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[4]_net_1 ));
    CFG4 #( .INIT(16'hFF10) )  \ahb_fsm_current_state_ns_0[0]  (.A(
        defSlaveSMNextState), .B(N_53), .C(N_63), .D(N_84), .Y(
        \ahb_fsm_current_state_ns[0] ));
    CFG4 #( .INIT(16'hEEEC) )  \ahb_fsm_current_state_ns_0[5]  (.A(
        \ahb_fsm_current_state[5]_net_1 ), .B(
        \ahb_fsm_current_state[4]_net_1 ), .C(N_53), .D(
        defSlaveSMNextState), .Y(\ahb_fsm_current_state_ns[5] ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[11]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[11])
        , .Y(\HADDR_6[11]_net_1 ));
    SLE \HWDATA_int[28]  (.D(eSRAM_eNVM_RW_0_DATAOUT[28]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[28]_net_1 ));
    CFG4 #( .INIT(16'hEEEC) )  \ahb_fsm_current_state_ns_0[2]  (.A(
        \ahb_fsm_current_state[2]_net_1 ), .B(
        \ahb_fsm_current_state[1]_net_1 ), .C(N_53), .D(
        defSlaveSMNextState), .Y(\ahb_fsm_current_state_ns[2] ));
    SLE \DATAOUT[29]  (.D(AHB_IF_0_BIF_1_HRDATA[29]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[29]));
    CFG4 #( .INIT(16'h0001) )  \ahb_fsm_current_state_ns_0_a2_0_1[0]  
        (.A(eSRAM_eNVM_RW_0_WRITE), .B(eSRAM_eNVM_RW_0_READ), .C(
        \ahb_fsm_current_state[2]_net_1 ), .D(
        \ahb_fsm_current_state[5]_net_1 ), .Y(N_52));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[12]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[12])
        , .Y(\HADDR_6[12]_net_1 ));
    SLE \DATAOUT[10]  (.D(AHB_IF_0_BIF_1_HRDATA[10]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[10]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[2]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[2]), 
        .Y(\HADDR_6[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[20]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[20])
        , .Y(\HADDR_6[20]_net_1 ));
    SLE \DATAOUT[6]  (.D(AHB_IF_0_BIF_1_HRDATA[6]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[6]));
    SLE \HWDATA_int[26]  (.D(eSRAM_eNVM_RW_0_DATAOUT[26]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[26]_net_1 ));
    SLE \HWDATA[27]  (.D(\HWDATA_int[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[27]));
    VCC VCC (.Y(VCC_net_1));
    SLE \HWDATA[8]  (.D(\HWDATA_int[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[8]));
    SLE \HWDATA_int[5]  (.D(eSRAM_eNVM_RW_0_DATAOUT[5]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[5]_net_1 ));
    SLE \HWDATA_int[11]  (.D(eSRAM_eNVM_RW_0_DATAOUT[11]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[11]_net_1 ));
    SLE \HADDR[22]  (.D(\HADDR_6[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[22]));
    SLE \HWDATA[18]  (.D(\HWDATA_int[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[18]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[31]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[31])
        , .Y(\HADDR_6[31]_net_1 ));
    SLE \HWDATA[15]  (.D(\HWDATA_int[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[15]));
    SLE \HWDATA[14]  (.D(\HWDATA_int[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[14]));
    SLE \HADDR[23]  (.D(\HADDR_6[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[23]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[25]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[25])
        , .Y(\HADDR_6[25]_net_1 ));
    SLE \DATAOUT[5]  (.D(AHB_IF_0_BIF_1_HRDATA[5]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[5]));
    SLE \HWDATA_int[13]  (.D(eSRAM_eNVM_RW_0_DATAOUT[13]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[13]_net_1 ));
    SLE \HWDATA[4]  (.D(\HWDATA_int[4]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[4]));
    SLE \DATAOUT[7]  (.D(AHB_IF_0_BIF_1_HRDATA[7]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[7]));
    SLE \HWDATA[7]  (.D(\HWDATA_int[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[7]));
    SLE \HWDATA[0]  (.D(\HWDATA_int[0]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[0]));
    SLE \HADDR[15]  (.D(\HADDR_6[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[15]));
    SLE \HWDATA[28]  (.D(\HWDATA_int[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[28]));
    SLE \HADDR[17]  (.D(\HADDR_6[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[17]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[16]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[16])
        , .Y(\HADDR_6[16]_net_1 ));
    SLE \HWDATA[11]  (.D(\HWDATA_int[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[11]));
    SLE \HWDATA[25]  (.D(\HWDATA_int[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[25]));
    SLE \DATAOUT[24]  (.D(AHB_IF_0_BIF_1_HRDATA[24]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[24]));
    SLE \HWDATA_int[10]  (.D(eSRAM_eNVM_RW_0_DATAOUT[10]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[10]_net_1 ));
    SLE \HADDR[11]  (.D(\HADDR_6[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[11]));
    SLE \DATAOUT[31]  (.D(AHB_IF_0_BIF_1_HRDATA[31]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[31]));
    SLE \HWDATA[24]  (.D(\HWDATA_int[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[24]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[24]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[24])
        , .Y(\HADDR_6[24]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \ahb_fsm_current_state_ns_0_o2[0]  (.A(
        \ahb_fsm_current_state[6]_net_1 ), .B(
        \ahb_fsm_current_state[3]_net_1 ), .Y(N_63));
    SLE \HWDATA_int[21]  (.D(eSRAM_eNVM_RW_0_DATAOUT[21]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[21]_net_1 ));
    SLE \HWDATA_int[14]  (.D(eSRAM_eNVM_RW_0_DATAOUT[14]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[14]_net_1 ));
    SLE \HADDR[16]  (.D(\HADDR_6[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[16]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[4]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[4]), 
        .Y(\HADDR_6[4]_net_1 ));
    SLE \HTRANS_1[1]  (.D(N_46), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(un1_N_5_mux_0_i_0), .ALn(eSRAM_eNVM_access_0_HPMS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(AHB_IF_0_BIF_1_HTRANS[1]));
    SLE \HWDATA_int[2]  (.D(eSRAM_eNVM_RW_0_DATAOUT[2]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[2]_net_1 ));
    SLE \HWDATA[31]  (.D(\HWDATA_int[31]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[31]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[21]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[21])
        , .Y(\HADDR_6[21]_net_1 ));
    CFG3 #( .INIT(8'h04) )  HWDATA_1_sqmuxa_0_a3_0_a2 (.A(N_53), .B(
        \ahb_fsm_current_state[2]_net_1 ), .C(defSlaveSMNextState), .Y(
        HWDATA_1_sqmuxa));
    SLE \HWDATA_int[6]  (.D(eSRAM_eNVM_RW_0_DATAOUT[6]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[6]_net_1 ));
    SLE \HWDATA[13]  (.D(\HWDATA_int[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[13]));
    CFG4 #( .INIT(16'hCCCE) )  VALID_RNO (.A(
        \ahb_fsm_current_state[6]_net_1 ), .B(
        \ahb_fsm_current_state[0]_net_1 ), .C(defSlaveSMNextState), .D(
        N_53), .Y(un18_N_5_mux_i_0));
    SLE \DATAOUT[15]  (.D(AHB_IF_0_BIF_1_HRDATA[15]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[15]));
    SLE \HWDATA_int[8]  (.D(eSRAM_eNVM_RW_0_DATAOUT[8]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[13]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[13])
        , .Y(\HADDR_6[13]_net_1 ));
    SLE \HADDR[31]  (.D(\HADDR_6[31]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[31]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[22]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[22])
        , .Y(\HADDR_6[22]_net_1 ));
    SLE \HWDATA_int[23]  (.D(eSRAM_eNVM_RW_0_DATAOUT[23]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[23]_net_1 ));
    CFG4 #( .INIT(16'hCCCE) )  HWRITE_RNO (.A(
        \ahb_fsm_current_state[2]_net_1 ), .B(N_115), .C(
        defSlaveSMNextState), .D(N_53), .Y(un1_N_5_mux_i_0));
    SLE \HWDATA[21]  (.D(\HWDATA_int[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[21]));
    CFG3 #( .INIT(8'h04) )  DATAOUT_1_sqmuxa_0_a3_0_a2 (.A(N_53), .B(
        \ahb_fsm_current_state[6]_net_1 ), .C(defSlaveSMNextState), .Y(
        DATAOUT_1_sqmuxa));
    SLE \DATAOUT[27]  (.D(AHB_IF_0_BIF_1_HRDATA[27]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[27]));
    SLE \HADDR[5]  (.D(\HADDR_6[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[5]));
    SLE \HADDR[25]  (.D(\HADDR_6[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[25]));
    SLE \HWDATA_int[31]  (.D(eSRAM_eNVM_RW_0_DATAOUT[31]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[31]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[6]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[6]), 
        .Y(\HADDR_6[6]_net_1 ));
    SLE \DATAOUT[4]  (.D(AHB_IF_0_BIF_1_HRDATA[4]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[4]));
    SLE \HWDATA[16]  (.D(\HWDATA_int[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[16]));
    SLE \HADDR[27]  (.D(\HADDR_6[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[27]));
    SLE \DATAOUT[11]  (.D(AHB_IF_0_BIF_1_HRDATA[11]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[11]));
    SLE \DATAOUT[12]  (.D(AHB_IF_0_BIF_1_HRDATA[12]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[12]));
    SLE \HWDATA_int[3]  (.D(eSRAM_eNVM_RW_0_DATAOUT[3]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[3]_net_1 ));
    SLE \HADDR[21]  (.D(\HADDR_6[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[21]));
    SLE \HWDATA_int[20]  (.D(eSRAM_eNVM_RW_0_DATAOUT[20]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[20]_net_1 ));
    SLE \HWDATA[1]  (.D(\HWDATA_int[1]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[1]));
    SLE HWRITE (.D(\ahb_fsm_current_state[1]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_N_5_mux_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWRITE));
    SLE \HADDR[26]  (.D(\HADDR_6[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[26]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[9]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[9]), 
        .Y(\HADDR_6[9]_net_1 ));
    SLE \HWDATA[23]  (.D(\HWDATA_int[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[23]));
    SLE \DATAOUT[9]  (.D(AHB_IF_0_BIF_1_HRDATA[9]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[9]));
    SLE \ahb_fsm_current_state[2]  (.D(\ahb_fsm_current_state_ns[2] ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[2]_net_1 ));
    SLE \HWDATA_int[24]  (.D(eSRAM_eNVM_RW_0_DATAOUT[24]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[24]_net_1 ));
    SLE \DATAOUT[13]  (.D(AHB_IF_0_BIF_1_HRDATA[13]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[13]));
    SLE \HWDATA_int[15]  (.D(eSRAM_eNVM_RW_0_DATAOUT[15]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[15]_net_1 ));
    SLE \HADDR[2]  (.D(\HADDR_6[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[2]));
    SLE \DATAOUT[20]  (.D(AHB_IF_0_BIF_1_HRDATA[20]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[20]));
    SLE \HWDATA_int[17]  (.D(eSRAM_eNVM_RW_0_DATAOUT[17]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[17]_net_1 ));
    SLE \HADDR[4]  (.D(\HADDR_6[4]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[4]));
    SLE \DATAOUT[18]  (.D(AHB_IF_0_BIF_1_HRDATA[18]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[18]));
    SLE \HWDATA[12]  (.D(\HWDATA_int[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[12]));
    SLE \HWDATA[26]  (.D(\HWDATA_int[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[26]));
    SLE \HWDATA_int[30]  (.D(eSRAM_eNVM_RW_0_DATAOUT[30]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[30]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[19]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[19])
        , .Y(\HADDR_6[19]_net_1 ));
    SLE \HWDATA_int[4]  (.D(eSRAM_eNVM_RW_0_DATAOUT[4]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[26]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[26])
        , .Y(\HADDR_6[26]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[18]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[18])
        , .Y(\HADDR_6[18]_net_1 ));
    SLE \HWDATA_int[12]  (.D(eSRAM_eNVM_RW_0_DATAOUT[12]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[12]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \ahb_fsm_current_state_ns_0_a2_0[0]  (
        .A(\ahb_fsm_current_state[3]_net_1 ), .B(
        \ahb_fsm_current_state[6]_net_1 ), .C(N_115), .D(N_52), .Y(
        N_84));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[17]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[17])
        , .Y(\HADDR_6[17]_net_1 ));
    SLE \HWDATA[10]  (.D(\HWDATA_int[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[10]));
    SLE \HADDR[14]  (.D(\HADDR_6[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[14]));
    SLE \HWDATA[19]  (.D(\HWDATA_int[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[19]));
    SLE \HADDR[10]  (.D(\HADDR_6[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[10]));
    CFG3 #( .INIT(8'h40) )  \ahb_fsm_current_state_ns_a3_0_a2[4]  (.A(
        eSRAM_eNVM_RW_0_WRITE), .B(\ahb_fsm_current_state[0]_net_1 ), 
        .C(eSRAM_eNVM_RW_0_READ), .Y(\ahb_fsm_current_state_ns[4] ));
    SLE \HWDATA_int[19]  (.D(eSRAM_eNVM_RW_0_DATAOUT[19]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[19]_net_1 ));
    SLE \HWDATA[22]  (.D(\HWDATA_int[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[22]));
    SLE \DATAOUT[16]  (.D(AHB_IF_0_BIF_1_HRDATA[16]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[16]));
    SLE \HWDATA[30]  (.D(\HWDATA_int[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[30]));
    SLE \HWDATA_int[25]  (.D(eSRAM_eNVM_RW_0_DATAOUT[25]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[25]_net_1 ));
    SLE \HWDATA[6]  (.D(\HWDATA_int[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[6]));
    SLE \HWDATA_int[27]  (.D(eSRAM_eNVM_RW_0_DATAOUT[27]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[27]_net_1 ));
    SLE \DATAOUT[8]  (.D(AHB_IF_0_BIF_1_HRDATA[8]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[8]));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[23]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[23])
        , .Y(\HADDR_6[23]_net_1 ));
    SLE \DATAOUT[19]  (.D(AHB_IF_0_BIF_1_HRDATA[19]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[19]));
    SLE \HADDR[30]  (.D(\HADDR_6[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[30]));
    SLE \HADDR[7]  (.D(\HADDR_6[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[7]));
    SLE \HWDATA[20]  (.D(\HWDATA_int[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[20]));
    SLE \HWDATA[29]  (.D(\HWDATA_int[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[29]));
    CFG4 #( .INIT(16'hEFE0) )  AHB_BUSY_RNO_0 (.A(eSRAM_eNVM_RW_0_READ)
        , .B(eSRAM_eNVM_RW_0_WRITE), .C(
        \ahb_fsm_current_state[0]_net_1 ), .D(N_63), .Y(N_106_i_0));
    CFG3 #( .INIT(8'hFB) )  un1_HADDR_0_sqmuxa_i_0_o2 (.A(N_53), .B(
        N_22), .C(defSlaveSMNextState), .Y(N_46));
    SLE VALID (.D(DATAOUT_1_sqmuxa), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un18_N_5_mux_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(AHB_IF_0_VALID)
        );
    CFG3 #( .INIT(8'h01) )  \HTRANS_1_RNO_0[1]  (.A(
        \ahb_fsm_current_state[1]_net_1 ), .B(
        \ahb_fsm_current_state[2]_net_1 ), .C(
        \ahb_fsm_current_state[4]_net_1 ), .Y(un1_m2_0_a2_0_0));
    CFG2 #( .INIT(4'hE) )  un1_ahb_fsm_current_state_4_0_o3_0_o2 (.A(
        \ahb_fsm_current_state[1]_net_1 ), .B(
        \ahb_fsm_current_state[4]_net_1 ), .Y(N_115));
    SLE \ahb_fsm_current_state[0]  (.D(\ahb_fsm_current_state_ns[0] ), 
        .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \HADDR_6[7]  (.A(
        \ahb_fsm_current_state[0]_net_1 ), .B(eSRAM_eNVM_RW_0_ADDR[7]), 
        .Y(\HADDR_6[7]_net_1 ));
    SLE \HADDR[24]  (.D(\HADDR_6[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[24]));
    SLE \HWDATA[9]  (.D(\HWDATA_int[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HWDATA_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HWDATA[9]));
    SLE \HWDATA_int[22]  (.D(eSRAM_eNVM_RW_0_DATAOUT[22]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_47_i_0), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\HWDATA_int[22]_net_1 ));
    SLE \HADDR[20]  (.D(\HADDR_6[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_101_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_BIF_1_HADDR[20]));
    SLE \DATAOUT[25]  (.D(AHB_IF_0_BIF_1_HRDATA[25]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(DATAOUT_1_sqmuxa), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        AHB_IF_0_DATAOUT[25]));
    SLE \ahb_fsm_current_state[6]  (.D(
        \ahb_fsm_current_state[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(HREADY_M_0_iv_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ahb_fsm_current_state[6]_net_1 ));
    
endmodule


module SPI_Master(
       state,
       eSRAM_eNVM_RW_0_ram_waddr,
       PRDATA_c,
       eSRAM_eNVM_RW_0_ram_wdata,
       PWRITE_c,
       eSRAM_eNVM_access_0_FIC_0_CLK,
       MISO_c,
       eSRAM_eNVM_access_0_HPMS_READY,
       CLKOUT_cl,
       CLKOUT_1,
       MOSI_1,
       ss_n_c,
       CS_c,
       MOSI_cl
    );
output [0:0] state;
input  [4:0] eSRAM_eNVM_RW_0_ram_waddr;
output [31:0] PRDATA_c;
input  [31:0] eSRAM_eNVM_RW_0_ram_wdata;
input  PWRITE_c;
input  eSRAM_eNVM_access_0_FIC_0_CLK;
input  MISO_c;
input  eSRAM_eNVM_access_0_HPMS_READY;
output CLKOUT_cl;
output CLKOUT_1;
output MOSI_1;
output ss_n_c;
output CS_c;
output MOSI_cl;

    wire PWRITE_c_i_0, \state_i_0[0] , \slv_select[0]_net_1 , 
        VCC_net_1, PWDATA_buf_0_sqmuxa, GND_net_1, 
        \slv_select[1]_net_1 , \slv_select[2]_net_1 , 
        \slv_select[3]_net_1 , \slv_select[4]_net_1 , 
        \PRDATA_buf[17]_net_1 , \PRDATA_buf[16]_net_1 , 
        PRDATA_buf_0_sqmuxa_1, \PRDATA_buf[18]_net_1 , 
        \PRDATA_buf[19]_net_1 , \PRDATA_buf[20]_net_1 , 
        \PRDATA_buf[21]_net_1 , \PRDATA_buf[22]_net_1 , 
        \PRDATA_buf[23]_net_1 , \PRDATA_buf[24]_net_1 , 
        \PRDATA_buf[25]_net_1 , \PRDATA_buf[26]_net_1 , 
        \PRDATA_buf[27]_net_1 , \PRDATA_buf[28]_net_1 , 
        \PRDATA_buf[29]_net_1 , \PRDATA_buf[30]_net_1 , 
        \PRDATA_buf[31]_net_1 , \PRDATA_buf[2]_net_1 , 
        \PRDATA_buf[1]_net_1 , \PRDATA_buf[3]_net_1 , 
        \PRDATA_buf[4]_net_1 , \PRDATA_buf[5]_net_1 , 
        \PRDATA_buf[6]_net_1 , \PRDATA_buf[7]_net_1 , 
        \PRDATA_buf[8]_net_1 , \PRDATA_buf[9]_net_1 , 
        \PRDATA_buf[10]_net_1 , \PRDATA_buf[11]_net_1 , 
        \PRDATA_buf[12]_net_1 , \PRDATA_buf[13]_net_1 , 
        \PRDATA_buf[14]_net_1 , \PRDATA_buf[15]_net_1 , 
        \PWDATA_buf[27]_net_1 , \PWDATA_buf_RNO[27]_net_1 , 
        un1_reset_inv_2_i_0_net_1, \PWDATA_buf[28]_net_1 , 
        \PWDATA_buf_RNO[28]_net_1 , \PWDATA_buf[29]_net_1 , 
        \PWDATA_buf_RNO[29]_net_1 , \PWDATA_buf[30]_net_1 , 
        \PWDATA_buf_RNO[30]_net_1 , \PWDATA_buf[31]_net_1 , 
        \PWDATA_buf_RNO[31]_net_1 , \PWDATA_buf[32]_net_1 , N_329_i_0, 
        \PWDATA_buf[33]_net_1 , N_317_i_0, \PWDATA_buf[34]_net_1 , 
        N_328_i_0, \PWDATA_buf[35]_net_1 , N_316_i_0, 
        \PWDATA_buf[36]_net_1 , N_201_i_0, \PWDATA_buf[37]_net_1 , 
        N_899, \PWDATA_buf[38]_net_1 , \PWDATA_buf_RNO[38]_net_1 , 
        \PWDATA_buf[39]_net_1 , N_877, \PRDATA_buf[0]_net_1 , 
        \PWDATA_buf[12]_net_1 , \PWDATA_buf_RNO[12]_net_1 , 
        \PWDATA_buf[13]_net_1 , \PWDATA_buf_RNO[13]_net_1 , 
        \PWDATA_buf[14]_net_1 , \PWDATA_buf_RNO[14]_net_1 , 
        \PWDATA_buf[15]_net_1 , \PWDATA_buf_RNO[15]_net_1 , 
        \PWDATA_buf[16]_net_1 , \PWDATA_buf_RNO[16]_net_1 , 
        \PWDATA_buf[17]_net_1 , \PWDATA_buf_RNO[17]_net_1 , 
        \PWDATA_buf[18]_net_1 , \PWDATA_buf_RNO[18]_net_1 , 
        \PWDATA_buf[19]_net_1 , \PWDATA_buf_RNO[19]_net_1 , 
        \PWDATA_buf[20]_net_1 , \PWDATA_buf_RNO[20]_net_1 , 
        \PWDATA_buf[21]_net_1 , \PWDATA_buf_RNO[21]_net_1 , 
        \PWDATA_buf[22]_net_1 , \PWDATA_buf_RNO[22]_net_1 , 
        \PWDATA_buf[23]_net_1 , \PWDATA_buf_RNO[23]_net_1 , 
        \PWDATA_buf[24]_net_1 , \PWDATA_buf_RNO[24]_net_1 , 
        \PWDATA_buf[25]_net_1 , \PWDATA_buf_RNO[25]_net_1 , 
        \PWDATA_buf[26]_net_1 , \PWDATA_buf_RNO[26]_net_1 , N_315_i_0, 
        \PWDATA_buf[0]_net_1 , N_670_i_0, \PWDATA_buf[1]_net_1 , 
        \PWDATA_buf_RNO[1]_net_1 , \PWDATA_buf[2]_net_1 , 
        \PWDATA_buf_RNO[2]_net_1 , \PWDATA_buf[3]_net_1 , 
        \PWDATA_buf_RNO[3]_net_1 , \PWDATA_buf[4]_net_1 , 
        \PWDATA_buf_RNO[4]_net_1 , \PWDATA_buf[5]_net_1 , 
        \PWDATA_buf_RNO[5]_net_1 , \PWDATA_buf[6]_net_1 , 
        \PWDATA_buf_RNO[6]_net_1 , \PWDATA_buf[7]_net_1 , 
        \PWDATA_buf_RNO[7]_net_1 , \PWDATA_buf[8]_net_1 , 
        \PWDATA_buf_RNO[8]_net_1 , \PWDATA_buf[9]_net_1 , 
        \PWDATA_buf_RNO[9]_net_1 , \PWDATA_buf[10]_net_1 , 
        \PWDATA_buf_RNO[10]_net_1 , \PWDATA_buf[11]_net_1 , 
        \PWDATA_buf_RNO[11]_net_1 , \count[31]_net_1 , 
        \count_0[31]_net_1 , \count[16]_net_1 , \count_0[16]_net_1 , 
        \count[17]_net_1 , \count_0[17]_net_1 , \count[18]_net_1 , 
        \count_0[18]_net_1 , \count[19]_net_1 , \count_0[19]_net_1 , 
        \count[20]_net_1 , \count_0[20]_net_1 , \count[21]_net_1 , 
        \count_0[21]_net_1 , \count[22]_net_1 , \count_0[22]_net_1 , 
        \count[23]_net_1 , \count_0[23]_net_1 , \count[24]_net_1 , 
        \count_0[24]_net_1 , \count[25]_net_1 , \count_0[25]_net_1 , 
        \count[26]_net_1 , \count_0[26]_net_1 , \count[27]_net_1 , 
        \count_0[27]_net_1 , \count[28]_net_1 , \count_0[28]_net_1 , 
        \count[29]_net_1 , \count_0[29]_net_1 , \count[30]_net_1 , 
        \count_0[30]_net_1 , \count[1]_net_1 , N_173_i_0, 
        \count[2]_net_1 , \count_0[2]_net_1 , \count[3]_net_1 , 
        \count_0[3]_net_1 , \count[4]_net_1 , N_179_i_0, 
        \count[5]_net_1 , N_326_i_0, \count[6]_net_1 , 
        \count_0[6]_net_1 , \count[7]_net_1 , \count_0[7]_net_1 , 
        \count[8]_net_1 , \count_0[8]_net_1 , \count[9]_net_1 , 
        \count_0[9]_net_1 , \count[10]_net_1 , \count_0[10]_net_1 , 
        \count[11]_net_1 , \count_0[11]_net_1 , \count[12]_net_1 , 
        \count_0[12]_net_1 , \count[13]_net_1 , \count_0[13]_net_1 , 
        \count[14]_net_1 , \count_0[14]_net_1 , \count[15]_net_1 , 
        \count_0[15]_net_1 , \count[0]_net_1 , \count_0[0]_net_1 , 
        CLKOUT_cl_1, CLKOUT_8_1_iv_i_0, continue_net_1, continue_4, 
        N_126_i_0, assert_data_net_1, N_327_i_0, \command[2]_net_1 , 
        \command[0]_net_1 , CS_6, N_324_i_0, un22_countlto6, 
        clk_toggles_5, un22_countlto5, clk_toggles_4, un22_countlto4, 
        clk_toggles_3, \clk_toggles[3]_net_1 , clk_toggles_2, 
        \clk_toggles[2]_net_1 , clk_toggles_1, \clk_toggles[1]_net_1 , 
        clk_toggles_0, \clk_toggles[0]_net_1 , clk_toggles, 
        un1_clk_toggles_1_cry_0, \clk_toggles_RNIKLQI_Y[0] , 
        un2_count_net_1, un1_clk_toggles_1_cry_1, 
        \clk_toggles_RNIVRNM_S[1] , un1_clk_toggles_1_cry_2, 
        \clk_toggles_RNIB3LQ_S[2] , un1_clk_toggles_1_cry_3, 
        \clk_toggles_RNIOBIU_S[3] , un1_clk_toggles_1_cry_4, 
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIKK8M1_S, un1_m1_e_0_0, 
        \clk_toggles_r_RNO_S[6] , un1_clk_toggles_1_cry_5, 
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIHUUD2_S, un1_count_s_0_73_FCO, 
        un1_count_cry_0_net_1, un1_count_cry_0_S, 
        un1_count_cry_1_net_1, un1_count_cry_1_S, 
        un1_count_cry_2_net_1, un1_count_cry_2_S, 
        un1_count_cry_3_net_1, un1_count_cry_3_S, 
        un1_count_cry_4_net_1, un1_count_cry_4_S, 
        un1_count_cry_5_net_1, un1_count_cry_5_S, 
        un1_count_cry_6_net_1, un1_count_cry_6_S, 
        un1_count_cry_7_net_1, un1_count_cry_7_S, 
        un1_count_cry_8_net_1, un1_count_cry_8_S, 
        un1_count_cry_9_net_1, un1_count_cry_9_S, 
        un1_count_cry_10_net_1, un1_count_cry_10_S, 
        un1_count_cry_11_net_1, un1_count_cry_11_S, 
        un1_count_cry_12_net_1, un1_count_cry_12_S, 
        un1_count_cry_13_net_1, un1_count_cry_13_S, 
        un1_count_cry_14_net_1, un1_count_cry_14_S, 
        un1_count_cry_15_net_1, un1_count_cry_15_S, 
        un1_count_cry_16_net_1, un1_count_cry_16_S, 
        un1_count_cry_17_net_1, un1_count_cry_17_S, 
        un1_count_cry_18_net_1, un1_count_cry_18_S, 
        un1_count_cry_19_net_1, un1_count_cry_19_S, 
        un1_count_cry_20_net_1, un1_count_cry_20_S, 
        un1_count_cry_21_net_1, un1_count_cry_21_S, 
        un1_count_cry_22_net_1, un1_count_cry_22_S, 
        un1_count_cry_23_net_1, un1_count_cry_23_S, 
        un1_count_cry_24_net_1, un1_count_cry_24_S, 
        un1_count_cry_25_net_1, un1_count_cry_25_S, 
        un1_count_cry_26_net_1, un1_count_cry_26_S, 
        un1_count_cry_27_net_1, un1_count_cry_27_S, 
        un1_count_cry_28_net_1, un1_count_cry_28_S, 
        un1_count_cry_29_net_1, un1_count_cry_29_S, un1_count_s_31_S, 
        un1_count_cry_30_net_1, un1_count_cry_30_S, N_509, N_477, 
        clk_toggles_0_sqmuxa_1, N_344, 
        PRDATA_buf_0_sqmuxa_1_0_a2_1_net_1, 
        continue_4_iv_0_a2_0_0_net_1, CLKOUT_8_1_iv_0_a2_0_0, 
        un2_count_23_net_1, un2_count_22_net_1, un2_count_21_net_1, 
        un2_count_20_net_1, un2_count_19_net_1, un2_count_18_net_1, 
        un2_count_17_net_1, un2_count_16_net_1, N_529, 
        CLKOUT_8_1_iv_0_o2_0_1_net_1, 
        clk_toggles_0_sqmuxa_1_0_a2_0_0_net_1, N_350, 
        CLKOUT_cl_1_u_0_a2_0, un2_count_29_net_1, un2_count_28_net_1, 
        CLKOUT_8_1_iv_0_a2_1_2_net_1, N_515, 
        continue_4_iv_0_a2_0_1_net_1, N_388, N_420_2, 
        CLKOUT_8_1_iv_0_a2_2_2_net_1, N_353, CLKOUT_cl_1_u_0_0_1_net_1, 
        un1_pwdata_5_645_i_m2_i_0, un1_pwdata_7_609_i_m2_i_0, 
        un1_pwdata_8_591_i_m2_i_0, un1_pwdata_6_627_i_m2_i_0, 
        un1_pwdata_4_663_i_m2_i_0, N_483, CLKOUT_8_1_iv_0_0_net_1;
    
    CFG4 #( .INIT(16'h0001) )  un2_count_20 (.A(\count[15]_net_1 ), .B(
        \count[14]_net_1 ), .C(\count[13]_net_1 ), .D(
        \count[12]_net_1 ), .Y(un2_count_20_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[21]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[21]), .B(\PWDATA_buf[20]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[21]_net_1 ));
    CFG4 #( .INIT(16'h557F) )  PRDATA_buf_0_sqmuxa_1_0_o2 (.A(
        un22_countlto6), .B(un22_countlto4), .C(N_350), .D(
        un22_countlto5), .Y(N_388));
    CFG2 #( .INIT(4'h2) )  \count_0[8]  (.A(un1_count_cry_8_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[8]_net_1 ));
    SLE \count[27]  (.D(\count_0[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[27]_net_1 ));
    SLE \state[0]  (.D(VCC_net_1), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(VCC_net_1), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(state[0]));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[25]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[25]), .B(\PWDATA_buf[24]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[25]_net_1 ));
    SLE \PRDATA_buf[2]  (.D(\PRDATA_buf[1]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[2]_net_1 ));
    SLE \count[25]  (.D(\count_0[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[25]_net_1 ));
    CFG2 #( .INIT(4'hD) )  CLKOUT_cl_1_u_0_o2 (.A(ss_n_c), .B(PWRITE_c)
        , .Y(N_344));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_20 (.A(VCC_net_1), .B(
        \count[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_19_net_1), .S(un1_count_cry_20_S), .Y(), .FCO(
        un1_count_cry_20_net_1));
    CFG3 #( .INIT(8'hB3) )  CS_6_0 (.A(continue_net_1), .B(state[0]), 
        .C(un2_count_net_1), .Y(CS_6));
    SLE \count[17]  (.D(\count_0[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[17]_net_1 ));
    SLE \PWDATA_buf[4]  (.D(\PWDATA_buf_RNO[4]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[4]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[20]  (.A(un1_count_cry_20_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[20]_net_1 ));
    SLE \count[15]  (.D(\count_0[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[15]_net_1 ));
    SLE \PWDATA_buf[34]  (.D(N_328_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[34]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[20]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[20]), .B(\PWDATA_buf[19]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[20]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[31]  (.A(un1_count_s_31_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[31]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[9]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[9]), .B(\PWDATA_buf[8]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[9]_net_1 ));
    CFG4 #( .INIT(16'hF870) )  \PWDATA_buf_RNO[39]  (.A(state[0]), .B(
        N_515), .C(\command[2]_net_1 ), .D(\PWDATA_buf[38]_net_1 ), .Y(
        N_877));
    SLE \PWDATA_buf[12]  (.D(\PWDATA_buf_RNO[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[12]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[3]  (.A(un1_count_cry_3_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[3]_net_1 ));
    ARI1 #( .INIT(20'h52FD0) )  \clk_toggles_RNIKLQI[0]  (.A(
        \clk_toggles[0]_net_1 ), .B(state[0]), .C(un2_count_net_1), .D(
        eSRAM_eNVM_access_0_HPMS_READY), .FCI(GND_net_1), .S(), .Y(
        \clk_toggles_RNIKLQI_Y[0] ), .FCO(un1_clk_toggles_1_cry_0));
    SLE \count[9]  (.D(\count_0[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[9]_net_1 ));
    SLE \PRDATA[5]  (.D(\PRDATA_buf[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[5]));
    SLE \PRDATA[30]  (.D(\PRDATA_buf[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[30]));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_27 (.A(VCC_net_1), .B(
        \count[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_26_net_1), .S(un1_count_cry_27_S), .Y(), .FCO(
        un1_count_cry_27_net_1));
    SLE \PWDATA_buf[33]  (.D(N_317_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[33]_net_1 ));
    SLE \PRDATA_buf[28]  (.D(\PRDATA_buf[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[28]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[21]  (.A(un1_count_cry_21_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[21]_net_1 ));
    CFG3 #( .INIT(8'h2A) )  \PWDATA_buf_RNO[0]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[0]), .B(state[0]), .C(N_515), .Y(
        N_670_i_0));
    SLE \PWDATA_buf[10]  (.D(\PWDATA_buf_RNO[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[10]_net_1 ));
    CFG4 #( .INIT(16'hCECC) )  CLKOUT_cl_1_u_0_0 (.A(un2_count_net_1), 
        .B(CLKOUT_cl_1_u_0_0_1_net_1), .C(un22_countlto5), .D(N_420_2), 
        .Y(CLKOUT_cl_1));
    SLE \PWDATA_buf[21]  (.D(\PWDATA_buf_RNO[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[21]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[4]  (.A(
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIKK8M1_S), .B(
        clk_toggles_0_sqmuxa_1), .Y(clk_toggles_3));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_9 (.A(VCC_net_1), .B(
        \count[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_8_net_1), .S(un1_count_cry_9_S), .Y(), .FCO(
        un1_count_cry_9_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[7]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[7]), .B(\PWDATA_buf[6]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_2 (.A(VCC_net_1), .B(
        \count[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_1_net_1), .S(un1_count_cry_2_S), .Y(), .FCO(
        un1_count_cry_2_net_1));
    SLE \slv_select[4]  (.D(eSRAM_eNVM_RW_0_ram_waddr[4]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\slv_select[4]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[27]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[27]), .B(\PWDATA_buf[26]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[27]_net_1 ));
    SLE \PRDATA_buf[5]  (.D(\PRDATA_buf[4]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[5]_net_1 ));
    SLE \PWDATA_buf[35]  (.D(N_316_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[35]_net_1 ));
    SLE \PRDATA[28]  (.D(\PRDATA_buf[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[28]));
    SLE \count[8]  (.D(\count_0[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[8]_net_1 ));
    SLE \command[2]  (.D(PWRITE_c), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .EN(PWDATA_buf_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \command[2]_net_1 ));
    CFG4 #( .INIT(16'hFCDC) )  \count_RNO[1]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(PWDATA_buf_0_sqmuxa), .C(
        un1_count_cry_1_S), .D(N_353), .Y(N_173_i_0));
    SLE \PWDATA_buf[39]  (.D(N_877), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[39]_net_1 ));
    CFG4 #( .INIT(16'hC088) )  continue_4_iv_0_0 (.A(continue_net_1), 
        .B(state[0]), .C(continue_4_iv_0_a2_0_1_net_1), .D(
        un2_count_net_1), .Y(continue_4));
    SLE \PWDATA_buf[5]  (.D(\PWDATA_buf_RNO[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[1]  (.A(
        \clk_toggles_RNIVRNM_S[1] ), .B(clk_toggles_0_sqmuxa_1), .Y(
        clk_toggles_0));
    SLE \slv_select[2]  (.D(eSRAM_eNVM_RW_0_ram_waddr[2]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\slv_select[2]_net_1 ));
    SLE \PRDATA[16]  (.D(\PRDATA_buf[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[16]));
    SLE \PRDATA[21]  (.D(\PRDATA_buf[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[21]));
    SLE \PRDATA[22]  (.D(\PRDATA_buf[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[22]));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_29 (.A(VCC_net_1), .B(
        \count[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_28_net_1), .S(un1_count_cry_29_S), .Y(), .FCO(
        un1_count_cry_29_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[2]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[2]), .B(\PWDATA_buf[1]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[2]_net_1 ));
    SLE \count[20]  (.D(\count_0[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[20]_net_1 ));
    CFG4 #( .INIT(16'h00F1) )  CLKOUT_8_1_iv_i (.A(
        CLKOUT_8_1_iv_0_a2_1_2_net_1), .B(CLKOUT_8_1_iv_0_a2_2_2_net_1)
        , .C(N_353), .D(CLKOUT_8_1_iv_0_0_net_1), .Y(CLKOUT_8_1_iv_i_0)
        );
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[19]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[19]), .B(\PWDATA_buf[18]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_4 (.A(VCC_net_1), .B(
        \count[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_3_net_1), .S(un1_count_cry_4_S), .Y(), .FCO(
        un1_count_cry_4_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_16 (.A(VCC_net_1), .B(
        \count[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_15_net_1), .S(un1_count_cry_16_S), .Y(), .FCO(
        un1_count_cry_16_net_1));
    SLE \PRDATA_buf[17]  (.D(\PRDATA_buf[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[17]_net_1 ));
    SLE \count[10]  (.D(\count_0[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[10]_net_1 ));
    SLE \PWDATA_buf[11]  (.D(\PWDATA_buf_RNO[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[11]_net_1 ));
    SLE \PWDATA_buf[24]  (.D(\PWDATA_buf_RNO[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[24]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[23]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[23]), .B(\PWDATA_buf[22]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[23]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_10 (.A(VCC_net_1), .B(
        \count[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_9_net_1), .S(un1_count_cry_10_S), .Y(), .FCO(
        un1_count_cry_10_net_1));
    SLE \count[5]  (.D(N_326_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \count[5]_net_1 ));
    SLE \command[0]  (.D(PWRITE_c_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\command[0]_net_1 ));
    SLE \PRDATA_buf[12]  (.D(\PRDATA_buf[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[12]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[1]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[1]), .B(\PWDATA_buf[0]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[1]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[16]  (.A(un1_count_cry_16_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[16]_net_1 ));
    CFG4 #( .INIT(16'h3133) )  \PWDATA_buf_RNO[34]  (.A(N_515), .B(
        un1_pwdata_6_627_i_m2_i_0), .C(\PWDATA_buf[33]_net_1 ), .D(
        state[0]), .Y(N_328_i_0));
    SLE \PWDATA_buf[23]  (.D(\PWDATA_buf_RNO[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[23]_net_1 ));
    SLE \PRDATA[9]  (.D(\PRDATA_buf[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[9]));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_17 (.A(VCC_net_1), .B(
        \count[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_16_net_1), .S(un1_count_cry_17_S), .Y(), .FCO(
        un1_count_cry_17_net_1));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h4) )  clk_toggles_0_sqmuxa_1_0_a2 (.A(state[0]), 
        .B(eSRAM_eNVM_access_0_HPMS_READY), .Y(PWDATA_buf_0_sqmuxa));
    SLE \PRDATA[25]  (.D(\PRDATA_buf[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[25]));
    CFG3 #( .INIT(8'h7F) )  continue_0_sqmuxa_i_o2 (.A(
        un2_count_28_net_1), .B(state[0]), .C(un2_count_29_net_1), .Y(
        N_353));
    CFG2 #( .INIT(4'h2) )  \count_0[12]  (.A(un1_count_cry_12_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[12]_net_1 ));
    SLE \PRDATA_buf[30]  (.D(\PRDATA_buf[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[30]_net_1 ));
    SLE \PRDATA_buf[10]  (.D(\PRDATA_buf[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[10]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_0 (.A(VCC_net_1), .B(
        \count[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_s_0_73_FCO), .S(un1_count_cry_0_S), .Y(), .FCO(
        un1_count_cry_0_net_1));
    SLE \PWDATA_buf[25]  (.D(\PWDATA_buf_RNO[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[25]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[28]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[28]), .B(\PWDATA_buf[27]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[28]_net_1 ));
    SLE \PWDATA_buf[8]  (.D(\PWDATA_buf_RNO[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[8]_net_1 ));
    CFG4 #( .INIT(16'h4044) )  CLKOUT_8_1_iv_0_a2 (.A(CLKOUT_1), .B(
        state[0]), .C(CLKOUT_8_1_iv_0_o2_0_1_net_1), .D(
        un2_count_net_1), .Y(N_483));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_1 (.A(VCC_net_1), .B(
        \count[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_0_net_1), .S(un1_count_cry_1_S), .Y(), .FCO(
        un1_count_cry_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \clk_toggles_r_RNO[6]  (.A(VCC_net_1), 
        .B(un22_countlto6), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_clk_toggles_1_cry_5), .S(\clk_toggles_r_RNO_S[6] ), .Y(), 
        .FCO());
    CFG4 #( .INIT(16'h8000) )  CLKOUT_8_1_iv_0_a2_1_2 (.A(CLKOUT_cl), 
        .B(CLKOUT_1), .C(N_509), .D(N_344), .Y(
        CLKOUT_8_1_iv_0_a2_1_2_net_1));
    SLE \PWDATA_buf[29]  (.D(\PWDATA_buf_RNO[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[29]_net_1 ));
    SLE \PWDATA_buf[38]  (.D(\PWDATA_buf_RNO[38]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[38]_net_1 ));
    SLE \PWDATA_buf[14]  (.D(\PWDATA_buf_RNO[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[14]_net_1 ));
    SLE \count[4]  (.D(N_179_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \count[4]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[26]  (.A(un1_count_cry_26_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[26]_net_1 ));
    SLE \PRDATA[18]  (.D(\PRDATA_buf[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[18]));
    SLE \count[22]  (.D(\count_0[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[22]_net_1 ));
    SLE MOSI_1_inst_1 (.D(\PWDATA_buf[39]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_126_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(MOSI_1));
    SLE CLKOUT_cl_inst_1 (.D(CLKOUT_cl_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        eSRAM_eNVM_access_0_HPMS_READY), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CLKOUT_cl));
    SLE \count[12]  (.D(\count_0[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[12]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  CLKOUT_8_1_iv_0_a2_0_0_0 (.A(
        un22_countlto4), .B(un22_countlto6), .C(CLKOUT_1), .D(state[0])
        , .Y(CLKOUT_8_1_iv_0_a2_0_0));
    CFG4 #( .INIT(16'hFEFC) )  un1_reset_inv_2_i_0 (.A(un2_count_net_1)
        , .B(N_477), .C(PWDATA_buf_0_sqmuxa), .D(un1_m1_e_0_0), .Y(
        un1_reset_inv_2_i_0_net_1));
    SLE \count[0]  (.D(\count_0[0]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[0]_net_1 ));
    CFG3 #( .INIT(8'h48) )  assert_data_RNO (.A(assert_data_net_1), .B(
        state[0]), .C(un2_count_net_1), .Y(N_327_i_0));
    SLE \slv_select[3]  (.D(eSRAM_eNVM_RW_0_ram_waddr[3]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\slv_select[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[22]  (.A(un1_count_cry_22_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[22]_net_1 ));
    SLE \PWDATA_buf[13]  (.D(\PWDATA_buf_RNO[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[13]_net_1 ));
    SLE \PRDATA_buf[26]  (.D(\PRDATA_buf[25]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[26]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \clk_toggles_RNIOBIU[3]  (.A(VCC_net_1)
        , .B(\clk_toggles[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_clk_toggles_1_cry_2), .S(\clk_toggles_RNIOBIU_S[3] ), 
        .Y(), .FCO(un1_clk_toggles_1_cry_3));
    CFG4 #( .INIT(16'h8000) )  un1_reset_inv_2_i_a2 (.A(PWRITE_c), .B(
        eSRAM_eNVM_access_0_HPMS_READY), .C(N_509), .D(un2_count_net_1)
        , .Y(N_477));
    CFG4 #( .INIT(16'h8000) )  un2_count_29 (.A(un2_count_23_net_1), 
        .B(un2_count_22_net_1), .C(un2_count_21_net_1), .D(
        un2_count_20_net_1), .Y(un2_count_29_net_1));
    CFG4 #( .INIT(16'hFFFE) )  PWDATA_buf_2_sqmuxa_0_o2 (.A(
        \clk_toggles[3]_net_1 ), .B(\clk_toggles[2]_net_1 ), .C(
        \clk_toggles[1]_net_1 ), .D(\clk_toggles[0]_net_1 ), .Y(N_350));
    CFG4 #( .INIT(16'hFCDC) )  \count_RNO[5]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(PWDATA_buf_0_sqmuxa), .C(
        un1_count_cry_5_S), .D(N_353), .Y(N_326_i_0));
    SLE \PRDATA_buf[6]  (.D(\PRDATA_buf[5]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_19 (.A(VCC_net_1), .B(
        \count[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_18_net_1), .S(un1_count_cry_19_S), .Y(), .FCO(
        un1_count_cry_19_net_1));
    CFG3 #( .INIT(8'h08) )  PRDATA_buf_0_sqmuxa_1_0_a2 (.A(
        PRDATA_buf_0_sqmuxa_1_0_a2_1_net_1), .B(N_388), .C(N_353), .Y(
        PRDATA_buf_0_sqmuxa_1));
    SLE \PRDATA_buf[3]  (.D(\PRDATA_buf[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[3]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[5]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[5]), .B(\PWDATA_buf[4]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[5]_net_1 ));
    SLE \PRDATA[7]  (.D(\PRDATA_buf[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[7]));
    SLE \PRDATA[11]  (.D(\PRDATA_buf[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[11]));
    SLE \PRDATA[12]  (.D(\PRDATA_buf[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[12]));
    SLE \PRDATA_buf[31]  (.D(\PRDATA_buf[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[31]_net_1 ));
    SLE \PRDATA_buf[11]  (.D(\PRDATA_buf[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[11]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[14]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[14]), .B(\PWDATA_buf[13]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[14]_net_1 ));
    SLE \PWDATA_buf[15]  (.D(\PWDATA_buf_RNO[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[15]_net_1 ));
    SLE \PRDATA[29]  (.D(\PRDATA_buf[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[29]));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_5 (.A(VCC_net_1), .B(
        \count[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_4_net_1), .S(un1_count_cry_5_S), .Y(), .FCO(
        un1_count_cry_5_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[17]  (.A(un1_count_cry_17_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[17]_net_1 ));
    SLE \PWDATA_buf[19]  (.D(\PWDATA_buf_RNO[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[19]_net_1 ));
    SLE \PRDATA[6]  (.D(\PRDATA_buf[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[6]));
    CFG4 #( .INIT(16'h0800) )  PWDATA_buf_2_sqmuxa_0_a2_0 (.A(
        un22_countlto4), .B(un22_countlto6), .C(un22_countlto5), .D(
        eSRAM_eNVM_access_0_HPMS_READY), .Y(N_529));
    CFG2 #( .INIT(4'h2) )  \count_0[18]  (.A(un1_count_cry_18_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[18]_net_1 ));
    SLE \PRDATA[24]  (.D(\PRDATA_buf[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[24]));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[26]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[26]), .B(\PWDATA_buf[25]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[26]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0001) )  un2_count_18 (.A(\count[23]_net_1 ), .B(
        \count[22]_net_1 ), .C(\count[21]_net_1 ), .D(
        \count[20]_net_1 ), .Y(un2_count_18_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[0]  (.A(un1_count_cry_0_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[0]_net_1 ));
    CFG4 #( .INIT(16'hFBBB) )  CLKOUT_cl_1_u_0_0_1 (.A(CLKOUT_cl), .B(
        state[0]), .C(CLKOUT_cl_1_u_0_a2_0), .D(un2_count_net_1), .Y(
        CLKOUT_cl_1_u_0_0_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_8 (.A(VCC_net_1), .B(
        \count[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_7_net_1), .S(un1_count_cry_8_S), .Y(), .FCO(
        un1_count_cry_8_net_1));
    SLE \PRDATA[15]  (.D(\PRDATA_buf[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[15]));
    CFG2 #( .INIT(4'h2) )  \count_0[27]  (.A(un1_count_cry_27_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[27]_net_1 ));
    SLE \PWDATA_buf[28]  (.D(\PWDATA_buf_RNO[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[28]_net_1 ));
    SLE \count[23]  (.D(\count_0[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[23]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[31]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[31]), .B(\PWDATA_buf[30]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[31]_net_1 ));
    SLE \PWDATA_buf[7]  (.D(\PWDATA_buf_RNO[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[7]_net_1 ));
    SLE \count[13]  (.D(\count_0[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[13]_net_1 ));
    CFG4 #( .INIT(16'h3133) )  \PWDATA_buf_RNO[35]  (.A(N_515), .B(
        un1_pwdata_7_609_i_m2_i_0), .C(\PWDATA_buf[34]_net_1 ), .D(
        state[0]), .Y(N_316_i_0));
    SLE \PRDATA_buf[14]  (.D(\PRDATA_buf[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[14]_net_1 ));
    SLE \PRDATA_buf[0]  (.D(MISO_c), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[28]  (.A(un1_count_cry_28_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[28]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un2_count_22 (.A(\count[7]_net_1 ), .B(
        \count[6]_net_1 ), .C(\count[3]_net_1 ), .D(\count[2]_net_1 ), 
        .Y(un2_count_22_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[22]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[22]), .B(\PWDATA_buf[21]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[22]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_28 (.A(VCC_net_1), .B(
        \count[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_27_net_1), .S(un1_count_cry_28_S), .Y(), .FCO(
        un1_count_cry_28_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[30]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[30]), .B(\PWDATA_buf[29]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[30]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_s_0_73 (.A(VCC_net_1), .B(
        eSRAM_eNVM_access_0_HPMS_READY), .C(GND_net_1), .D(GND_net_1), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(un1_count_s_0_73_FCO));
    SLE \PWDATA_buf[6]  (.D(\PWDATA_buf_RNO[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[6]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[13]  (.A(un1_count_cry_13_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[13]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  CLKOUT_8_1_iv_0_a2_2_3 (.A(ss_n_c), .B(
        N_350), .C(PWRITE_c), .D(assert_data_net_1), .Y(N_420_2));
    SLE \PRDATA_buf[13]  (.D(\PRDATA_buf[12]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \clk_toggles_RNIB3LQ[2]  (.A(VCC_net_1)
        , .B(\clk_toggles[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_clk_toggles_1_cry_1), .S(\clk_toggles_RNIB3LQ_S[2] ), 
        .Y(), .FCO(un1_clk_toggles_1_cry_2));
    SLE continue (.D(continue_4), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(eSRAM_eNVM_access_0_HPMS_READY), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(continue_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_s_31 (.A(VCC_net_1), .B(
        \count[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_30_net_1), .S(un1_count_s_31_S), .Y(), .FCO());
    SLE \slv_select[0]  (.D(eSRAM_eNVM_RW_0_ram_waddr[0]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\slv_select[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[14]  (.A(un1_count_cry_14_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[14]_net_1 ));
    SLE \PWDATA_buf[1]  (.D(\PWDATA_buf_RNO[1]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[1]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  PRDATA_buf_0_sqmuxa_1_0_a2_1 (.A(
        assert_data_net_1), .B(PWRITE_c), .C(
        eSRAM_eNVM_access_0_HPMS_READY), .D(ss_n_c), .Y(
        PRDATA_buf_0_sqmuxa_1_0_a2_1_net_1));
    SLE \PWDATA_buf[9]  (.D(\PWDATA_buf_RNO[9]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[9]_net_1 ));
    SLE \PRDATA_buf[15]  (.D(\PRDATA_buf[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[15]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[9]  (.A(un1_count_cry_9_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[9]_net_1 ));
    CFG4 #( .INIT(16'hF870) )  \PWDATA_buf_RNO[37]  (.A(state[0]), .B(
        N_515), .C(\command[0]_net_1 ), .D(\PWDATA_buf[36]_net_1 ), .Y(
        N_899));
    SLE \PWDATA_buf[36]  (.D(N_201_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[36]_net_1 ));
    SLE \PWDATA_buf[18]  (.D(\PWDATA_buf_RNO[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[18]_net_1 ));
    SLE \count[1]  (.D(N_173_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \count[1]_net_1 ));
    CFG4 #( .INIT(16'h04CC) )  CLKOUT_cl_1_u_0_a2_1 (.A(un22_countlto4)
        , .B(assert_data_net_1), .C(un22_countlto5), .D(un22_countlto6)
        , .Y(N_509));
    SLE \slv_select[1]  (.D(eSRAM_eNVM_RW_0_ram_waddr[1]), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PWDATA_buf_0_sqmuxa), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\slv_select[1]_net_1 ));
    SLE \PRDATA[19]  (.D(\PRDATA_buf[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[19]));
    SLE \PRDATA_buf[19]  (.D(\PRDATA_buf[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[19]_net_1 ));
    SLE \PWDATA_buf[0]  (.D(N_670_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[0]_net_1 ));
    SLE \count[3]  (.D(\count_0[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[3]_net_1 ));
    SLE \clk_toggles[2]  (.D(clk_toggles_1), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clk_toggles[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[23]  (.A(un1_count_cry_23_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[23]_net_1 ));
    SLE \count[29]  (.D(\count_0[29]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[29]_net_1 ));
    CFG4 #( .INIT(16'hFFE0) )  CLKOUT_8_1_iv_0_0 (.A(PWRITE_c), .B(
        N_350), .C(CLKOUT_8_1_iv_0_a2_0_0), .D(N_483), .Y(
        CLKOUT_8_1_iv_0_0_net_1));
    CFG1 #( .INIT(2'h1) )  \command_RNO[0]  (.A(PWRITE_c), .Y(
        PWRITE_c_i_0));
    SLE \count[19]  (.D(\count_0[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[19]_net_1 ));
    CFG2 #( .INIT(4'h4) )  continue_RNI7VVF (.A(N_353), .B(
        continue_net_1), .Y(N_315_i_0));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[11]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[11]), .B(\PWDATA_buf[10]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[11]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  clk_toggles_0_sqmuxa_1_0 (.A(N_529), .B(
        clk_toggles_0_sqmuxa_1_0_a2_0_0_net_1), .C(un2_count_net_1), 
        .D(PWDATA_buf_0_sqmuxa), .Y(clk_toggles_0_sqmuxa_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_22 (.A(VCC_net_1), .B(
        \count[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_21_net_1), .S(un1_count_cry_22_S), .Y(), .FCO(
        un1_count_cry_22_net_1));
    SLE \PRDATA[14]  (.D(\PRDATA_buf[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[14]));
    CFG1 #( .INIT(2'h1) )  ss_n_RNO (.A(state[0]), .Y(\state_i_0[0] ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[15]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[15]), .B(\PWDATA_buf[14]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[15]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[24]  (.A(un1_count_cry_24_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[24]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_23 (.A(VCC_net_1), .B(
        \count[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_22_net_1), .S(un1_count_cry_23_S), .Y(), .FCO(
        un1_count_cry_23_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[10]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[10]), .B(\PWDATA_buf[9]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[10]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[2]  (.A(
        \clk_toggles_RNIB3LQ_S[2] ), .B(clk_toggles_0_sqmuxa_1), .Y(
        clk_toggles_1));
    SLE \clk_toggles[0]  (.D(clk_toggles), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clk_toggles[0]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un2_count_16 (.A(\count[31]_net_1 ), .B(
        \count[30]_net_1 ), .C(\count[29]_net_1 ), .D(
        \count[28]_net_1 ), .Y(un2_count_16_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[4]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[4]), .B(\PWDATA_buf[3]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  MOSI_1_RNO (.A(N_353), .B(N_515), .Y(
        N_126_i_0));
    CFG2 #( .INIT(4'h2) )  \count_0[2]  (.A(un1_count_cry_2_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[2]_net_1 ));
    SLE \PRDATA[0]  (.D(\PRDATA_buf[0]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[0]));
    SLE \PRDATA[31]  (.D(\PRDATA_buf[31]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[31]));
    SLE \clk_toggles[1]  (.D(clk_toggles_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clk_toggles[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_6 (.A(VCC_net_1), .B(
        \count[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_5_net_1), .S(un1_count_cry_6_S), .Y(), .FCO(
        un1_count_cry_6_net_1));
    SLE \PRDATA_buf[27]  (.D(\PRDATA_buf[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[27]_net_1 ));
    CFG4 #( .INIT(16'h3133) )  \PWDATA_buf_RNO[33]  (.A(N_515), .B(
        un1_pwdata_5_645_i_m2_i_0), .C(\PWDATA_buf[32]_net_1 ), .D(
        state[0]), .Y(N_317_i_0));
    CFG2 #( .INIT(4'h8) )  un2_count (.A(un2_count_28_net_1), .B(
        un2_count_29_net_1), .Y(un2_count_net_1));
    SLE \PRDATA_buf[4]  (.D(\PRDATA_buf[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_18 (.A(VCC_net_1), .B(
        \count[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_17_net_1), .S(un1_count_cry_18_S), .Y(), .FCO(
        un1_count_cry_18_net_1));
    SLE \PRDATA[4]  (.D(\PRDATA_buf[4]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[4]));
    SLE CS (.D(CS_6), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        VCC_net_1), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CS_c));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_25 (.A(VCC_net_1), .B(
        \count[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_24_net_1), .S(un1_count_cry_25_S), .Y(), .FCO(
        un1_count_cry_25_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[17]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[17]), .B(\PWDATA_buf[16]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[17]_net_1 ));
    SLE \PRDATA_buf[22]  (.D(\PRDATA_buf[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[22]_net_1 ));
    CFG4 #( .INIT(16'h0533) )  \PWDATA_buf_RNO_0[32]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[0]), .B(\slv_select[0]_net_1 ), .C(
        N_515), .D(state[0]), .Y(un1_pwdata_4_663_i_m2_i_0));
    CFG4 #( .INIT(16'hFCDC) )  \count_RNO[4]  (.A(
        eSRAM_eNVM_access_0_HPMS_READY), .B(PWDATA_buf_0_sqmuxa), .C(
        un1_count_cry_4_S), .D(N_353), .Y(N_179_i_0));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[5]  (.A(
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIHUUD2_S), .B(
        clk_toggles_0_sqmuxa_1), .Y(clk_toggles_4));
    ARI1 #( .INIT(20'h4AA00) )  \clk_toggles_RNIVRNM[1]  (.A(VCC_net_1)
        , .B(\clk_toggles[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_clk_toggles_1_cry_0), .S(\clk_toggles_RNIVRNM_S[1] ), 
        .Y(), .FCO(un1_clk_toggles_1_cry_1));
    CFG2 #( .INIT(4'h2) )  PWDATA_buf_2_sqmuxa_0_a2_0_1 (.A(N_529), .B(
        N_350), .Y(un1_m1_e_0_0));
    SLE \PRDATA[20]  (.D(\PRDATA_buf[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[20]));
    SLE \PRDATA_buf[9]  (.D(\PRDATA_buf[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[9]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un2_count_21 (.A(\count[11]_net_1 ), .B(
        \count[10]_net_1 ), .C(\count[9]_net_1 ), .D(\count[8]_net_1 ), 
        .Y(un2_count_21_net_1));
    SLE \PWDATA_buf[26]  (.D(\PWDATA_buf_RNO[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[26]_net_1 ));
    CFG3 #( .INIT(8'hF7) )  \PWDATA_buf_RNO[38]  (.A(state[0]), .B(
        N_515), .C(\PWDATA_buf[37]_net_1 ), .Y(
        \PWDATA_buf_RNO[38]_net_1 ));
    SLE \PRDATA[2]  (.D(\PRDATA_buf[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[2]));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[29]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[29]), .B(\PWDATA_buf[28]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[29]_net_1 ));
    SLE CLKOUT_1_inst_1 (.D(CLKOUT_8_1_iv_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(
        eSRAM_eNVM_access_0_HPMS_READY), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CLKOUT_1));
    SLE \PRDATA_buf[20]  (.D(\PRDATA_buf[19]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[20]_net_1 ));
    SLE \PRDATA_buf[18]  (.D(\PRDATA_buf[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[18]_net_1 ));
    CFG3 #( .INIT(8'h40) )  continue_4_iv_0_a2_0_0 (.A(continue_net_1), 
        .B(un22_countlto4), .C(un22_countlto6), .Y(
        continue_4_iv_0_a2_0_0_net_1));
    ARI1 #( .INIT(20'h56AAA) )  PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIKK8M1 
        (.A(state[0]), .B(un22_countlto4), .C(un1_m1_e_0_0), .D(
        un2_count_net_1), .FCI(un1_clk_toggles_1_cry_3), .S(
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIKK8M1_S), .Y(), .FCO(
        un1_clk_toggles_1_cry_4));
    CFG2 #( .INIT(4'h2) )  \count_0[7]  (.A(un1_count_cry_7_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[7]_net_1 ));
    CFG4 #( .INIT(16'hBF3F) )  CLKOUT_8_1_iv_0_o2_0_1 (.A(
        un22_countlto6), .B(assert_data_net_1), .C(N_344), .D(
        un22_countlto5), .Y(CLKOUT_8_1_iv_0_o2_0_1_net_1));
    SLE \PRDATA[23]  (.D(\PRDATA_buf[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[23]));
    SLE \PRDATA[8]  (.D(\PRDATA_buf[8]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[8]));
    ARI1 #( .INIT(20'h56AAA) )  PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIHUUD2 
        (.A(state[0]), .B(un22_countlto5), .C(un1_m1_e_0_0), .D(
        un2_count_net_1), .FCI(un1_clk_toggles_1_cry_4), .S(
        PWDATA_buf_2_sqmuxa_0_a2_0_1_RNIHUUD2_S), .Y(), .FCO(
        un1_clk_toggles_1_cry_5));
    CFG4 #( .INIT(16'h0533) )  \PWDATA_buf_RNO_0[36]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[4]), .B(\slv_select[4]_net_1 ), .C(
        N_515), .D(state[0]), .Y(un1_pwdata_8_591_i_m2_i_0));
    SLE \clk_toggles[4]  (.D(clk_toggles_3), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(un22_countlto4));
    SLE \PRDATA_buf[7]  (.D(\PRDATA_buf[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_12 (.A(VCC_net_1), .B(
        \count[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_11_net_1), .S(un1_count_cry_12_S), .Y(), .FCO(
        un1_count_cry_12_net_1));
    CFG4 #( .INIT(16'h8000) )  un2_count_28 (.A(un2_count_19_net_1), 
        .B(un2_count_18_net_1), .C(un2_count_17_net_1), .D(
        un2_count_16_net_1), .Y(un2_count_28_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[13]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[13]), .B(\PWDATA_buf[12]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_24 (.A(VCC_net_1), .B(
        \count[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_23_net_1), .S(un1_count_cry_24_S), .Y(), .FCO(
        un1_count_cry_24_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[19]  (.A(un1_count_cry_19_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_30 (.A(VCC_net_1), .B(
        \count[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_29_net_1), .S(un1_count_cry_30_S), .Y(), .FCO(
        un1_count_cry_30_net_1));
    SLE \PRDATA_buf[1]  (.D(\PRDATA_buf[0]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_13 (.A(VCC_net_1), .B(
        \count[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_12_net_1), .S(un1_count_cry_13_S), .Y(), .FCO(
        un1_count_cry_13_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[15]  (.A(un1_count_cry_15_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[15]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[6]  (.A(un1_count_cry_6_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[6]_net_1 ));
    SLE \PWDATA_buf[16]  (.D(\PWDATA_buf_RNO[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[16]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  clk_toggles_0_sqmuxa_1_0_a2_0_0 (.A(
        \clk_toggles[3]_net_1 ), .B(\clk_toggles[2]_net_1 ), .C(
        \clk_toggles[1]_net_1 ), .D(\clk_toggles[0]_net_1 ), .Y(
        clk_toggles_0_sqmuxa_1_0_a2_0_0_net_1));
    SLE \PRDATA_buf[21]  (.D(\PRDATA_buf[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[21]_net_1 ));
    SLE \count[31]  (.D(\count_0[31]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[31]_net_1 ));
    SLE \count[28]  (.D(\count_0[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[28]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_21 (.A(VCC_net_1), .B(
        \count[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_20_net_1), .S(un1_count_cry_21_S), .Y(), .FCO(
        un1_count_cry_21_net_1));
    SLE \count[18]  (.D(\count_0[18]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[18]_net_1 ));
    SLE \PRDATA[27]  (.D(\PRDATA_buf[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[27]));
    SLE \PRDATA[1]  (.D(\PRDATA_buf[1]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[1]));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[18]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[18]), .B(\PWDATA_buf[17]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[18]_net_1 ));
    SLE \PRDATA_buf[8]  (.D(\PRDATA_buf[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[8]_net_1 ));
    SLE \PRDATA[3]  (.D(\PRDATA_buf[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[3]));
    SLE \count[7]  (.D(\count_0[7]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[7]_net_1 ));
    CFG4 #( .INIT(16'h3133) )  \PWDATA_buf_RNO[36]  (.A(N_515), .B(
        un1_pwdata_8_591_i_m2_i_0), .C(\PWDATA_buf[35]_net_1 ), .D(
        state[0]), .Y(N_201_i_0));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_15 (.A(VCC_net_1), .B(
        \count[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_14_net_1), .S(un1_count_cry_15_S), .Y(), .FCO(
        un1_count_cry_15_net_1));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[3]  (.A(
        \clk_toggles_RNIOBIU_S[3] ), .B(clk_toggles_0_sqmuxa_1), .Y(
        clk_toggles_2));
    CFG2 #( .INIT(4'h2) )  \count_0[29]  (.A(un1_count_cry_29_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[29]_net_1 ));
    SLE \PWDATA_buf[37]  (.D(N_899), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[37]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_3 (.A(VCC_net_1), .B(
        \count[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_2_net_1), .S(un1_count_cry_3_S), .Y(), .FCO(
        un1_count_cry_3_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[25]  (.A(un1_count_cry_25_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[25]_net_1 ));
    CFG3 #( .INIT(8'h04) )  continue_4_iv_0_a2_0_1 (.A(un22_countlto5), 
        .B(continue_4_iv_0_a2_0_0_net_1), .C(N_350), .Y(
        continue_4_iv_0_a2_0_1_net_1));
    CFG4 #( .INIT(16'h0080) )  un2_count_23 (.A(\count[5]_net_1 ), .B(
        \count[4]_net_1 ), .C(\count[1]_net_1 ), .D(\count[0]_net_1 ), 
        .Y(un2_count_23_net_1));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[3]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[3]), .B(\PWDATA_buf[2]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[3]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[8]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[8]), .B(\PWDATA_buf[7]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[8]_net_1 ));
    SLE \PRDATA[10]  (.D(\PRDATA_buf[10]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[10]));
    SLE \count[6]  (.D(\count_0[6]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[6]_net_1 ));
    SLE \PWDATA_buf[3]  (.D(\PWDATA_buf_RNO[3]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[3]_net_1 ));
    SLE \PWDATA_buf[2]  (.D(\PWDATA_buf_RNO[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[2]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[24]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[24]), .B(\PWDATA_buf[23]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[24]_net_1 ));
    SLE \PWDATA_buf[32]  (.D(N_329_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[32]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[6]  (.A(
        \clk_toggles_r_RNO_S[6] ), .B(clk_toggles_0_sqmuxa_1), .Y(
        clk_toggles_5));
    CFG4 #( .INIT(16'h0533) )  \PWDATA_buf_RNO_0[35]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[3]), .B(\slv_select[3]_net_1 ), .C(
        N_515), .D(state[0]), .Y(un1_pwdata_7_609_i_m2_i_0));
    CFG4 #( .INIT(16'h3133) )  \PWDATA_buf_RNO[32]  (.A(N_515), .B(
        un1_pwdata_4_663_i_m2_i_0), .C(\PWDATA_buf[31]_net_1 ), .D(
        state[0]), .Y(N_329_i_0));
    SLE \PRDATA_buf[24]  (.D(\PRDATA_buf[23]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[24]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  CLKOUT_8_1_iv_0_a2_2_2 (.A(CLKOUT_cl), 
        .B(un22_countlto5), .C(N_420_2), .D(CLKOUT_1), .Y(
        CLKOUT_8_1_iv_0_a2_2_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_7 (.A(VCC_net_1), .B(
        \count[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_6_net_1), .S(un1_count_cry_7_S), .Y(), .FCO(
        un1_count_cry_7_net_1));
    SLE \PWDATA_buf[30]  (.D(\PWDATA_buf_RNO[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[30]_net_1 ));
    SLE \PRDATA[13]  (.D(\PRDATA_buf[13]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[13]));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_14 (.A(VCC_net_1), .B(
        \count[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_13_net_1), .S(un1_count_cry_14_S), .Y(), .FCO(
        un1_count_cry_14_net_1));
    SLE \count[26]  (.D(\count_0[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[26]_net_1 ));
    SLE \PRDATA_buf[23]  (.D(\PRDATA_buf[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[23]_net_1 ));
    SLE \count[16]  (.D(\count_0[16]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[16]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un2_count_17 (.A(\count[27]_net_1 ), .B(
        \count[26]_net_1 ), .C(\count[25]_net_1 ), .D(
        \count[24]_net_1 ), .Y(un2_count_17_net_1));
    SLE \PRDATA_buf[16]  (.D(\PRDATA_buf[15]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[16]_net_1 ));
    SLE \count[2]  (.D(\count_0[2]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[2]_net_1 ));
    SLE \clk_toggles[5]  (.D(clk_toggles_4), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(un22_countlto5));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[16]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[16]), .B(\PWDATA_buf[15]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[16]_net_1 ));
    SLE \PRDATA_buf[25]  (.D(\PRDATA_buf[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[25]_net_1 ));
    SLE \clk_toggles[3]  (.D(clk_toggles_2), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clk_toggles[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_11 (.A(VCC_net_1), .B(
        \count[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_10_net_1), .S(un1_count_cry_11_S), .Y(), .FCO(
        un1_count_cry_11_net_1));
    SLE \PWDATA_buf[27]  (.D(\PWDATA_buf_RNO[27]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[27]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \clk_toggles_r[0]  (.A(
        \clk_toggles_RNIKLQI_Y[0] ), .B(clk_toggles_0_sqmuxa_1), .Y(
        clk_toggles));
    SLE \PRDATA_buf[29]  (.D(\PRDATA_buf[28]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(PRDATA_buf_0_sqmuxa_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PRDATA_buf[29]_net_1 ));
    SLE \count[21]  (.D(\count_0[21]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[21]_net_1 ));
    CFG2 #( .INIT(4'h8) )  un1_reset_inv_2_i_a2_1 (.A(N_509), .B(
        PWRITE_c), .Y(N_515));
    SLE MOSI_cl_inst_1 (.D(N_324_i_0), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(MOSI_cl));
    SLE \count[11]  (.D(\count_0[11]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[11]_net_1 ));
    SLE \PRDATA[17]  (.D(\PRDATA_buf[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[17]));
    CFG2 #( .INIT(4'h8) )  CLKOUT_cl_1_u_0_a2_0_0 (.A(N_344), .B(N_509)
        , .Y(CLKOUT_cl_1_u_0_a2_0));
    SLE \PWDATA_buf[31]  (.D(\PWDATA_buf_RNO[31]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[31]_net_1 ));
    SLE \clk_toggles[6]  (.D(clk_toggles_5), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(un22_countlto6));
    CFG4 #( .INIT(16'h0533) )  \PWDATA_buf_RNO_0[34]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[2]), .B(\slv_select[2]_net_1 ), .C(
        N_515), .D(state[0]), .Y(un1_pwdata_6_627_i_m2_i_0));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[12]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[12]), .B(\PWDATA_buf[11]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[12]_net_1 ));
    SLE \count[24]  (.D(\count_0[24]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[24]_net_1 ));
    SLE ss_n (.D(\state_i_0[0] ), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK), 
        .EN(VCC_net_1), .ALn(eSRAM_eNVM_access_0_HPMS_READY), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(ss_n_c));
    SLE \count[14]  (.D(\count_0[14]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[14]_net_1 ));
    SLE \PWDATA_buf[22]  (.D(\PWDATA_buf_RNO[22]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[22]_net_1 ));
    SLE \PRDATA[26]  (.D(\PRDATA_buf[26]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(N_315_i_0), .ALn(
        eSRAM_eNVM_access_0_HPMS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_c[26]));
    CFG2 #( .INIT(4'h2) )  \count_0[10]  (.A(un1_count_cry_10_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[10]_net_1 ));
    CFG4 #( .INIT(16'h0533) )  \PWDATA_buf_RNO_0[33]  (.A(
        eSRAM_eNVM_RW_0_ram_waddr[1]), .B(\slv_select[1]_net_1 ), .C(
        N_515), .D(state[0]), .Y(un1_pwdata_5_645_i_m2_i_0));
    SLE \count[30]  (.D(\count_0[30]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(VCC_net_1), .ALn(VCC_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count[30]_net_1 ));
    CFG4 #( .INIT(16'hC888) )  MOSI_cl_RNO (.A(MOSI_cl), .B(state[0]), 
        .C(N_515), .D(un2_count_net_1), .Y(N_324_i_0));
    CFG4 #( .INIT(16'h0001) )  un2_count_19 (.A(\count[19]_net_1 ), .B(
        \count[18]_net_1 ), .C(\count[17]_net_1 ), .D(
        \count[16]_net_1 ), .Y(un2_count_19_net_1));
    SLE \PWDATA_buf[20]  (.D(\PWDATA_buf_RNO[20]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[20]_net_1 ));
    SLE assert_data (.D(N_327_i_0), .CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .EN(eSRAM_eNVM_access_0_HPMS_READY), .ALn(VCC_net_1), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(assert_data_net_1));
    CFG2 #( .INIT(4'h2) )  \count_0[30]  (.A(un1_count_cry_30_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[30]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_count_cry_26 (.A(VCC_net_1), .B(
        \count[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_count_cry_25_net_1), .S(un1_count_cry_26_S), .Y(), .FCO(
        un1_count_cry_26_net_1));
    SLE \PWDATA_buf[17]  (.D(\PWDATA_buf_RNO[17]_net_1 ), .CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .EN(un1_reset_inv_2_i_0_net_1), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\PWDATA_buf[17]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \count_0[11]  (.A(un1_count_cry_11_S), .B(
        PWDATA_buf_0_sqmuxa), .Y(\count_0[11]_net_1 ));
    CFG4 #( .INIT(16'hCAAA) )  \PWDATA_buf_RNO[6]  (.A(
        eSRAM_eNVM_RW_0_ram_wdata[6]), .B(\PWDATA_buf[5]_net_1 ), .C(
        N_515), .D(state[0]), .Y(\PWDATA_buf_RNO[6]_net_1 ));
    
endmodule


module eSRAM_eNVM_access_top(
       PRDATA,
       RD,
       DEVRST_N,
       FAB_RESET_N,
       MISO,
       PWRITE,
       start_esram,
       CLKOUT,
       CS,
       MOSI,
       ss_n
    );
output [31:0] PRDATA;
output [7:0] RD;
input  DEVRST_N;
input  FAB_RESET_N;
input  MISO;
input  PWRITE;
input  start_esram;
output CLKOUT;
output CS;
output MOSI;
output ss_n;

    wire eSRAM_eNVM_access_0_FIC_0_CLK, eSRAM_eNVM_access_0_HPMS_READY, 
        eSRAM_eNVM_RW_0_READ, eSRAM_eNVM_RW_0_WRITE, 
        \eSRAM_eNVM_RW_0_ADDR[2] , \eSRAM_eNVM_RW_0_DATAOUT[0] , 
        GND_net_1, VCC_net_1, \AHB_IF_0_DATAOUT[0] , 
        \AHB_IF_0_DATAOUT[1] , \AHB_IF_0_DATAOUT[2] , 
        \AHB_IF_0_DATAOUT[3] , \AHB_IF_0_DATAOUT[4] , 
        \AHB_IF_0_DATAOUT[5] , \AHB_IF_0_DATAOUT[6] , 
        \AHB_IF_0_DATAOUT[7] , \AHB_IF_0_DATAOUT[8] , 
        \AHB_IF_0_DATAOUT[9] , \AHB_IF_0_DATAOUT[10] , 
        \AHB_IF_0_DATAOUT[11] , \AHB_IF_0_DATAOUT[12] , 
        \AHB_IF_0_DATAOUT[13] , \AHB_IF_0_DATAOUT[14] , 
        \AHB_IF_0_DATAOUT[15] , \AHB_IF_0_DATAOUT[16] , 
        \AHB_IF_0_DATAOUT[17] , \AHB_IF_0_DATAOUT[18] , 
        \AHB_IF_0_DATAOUT[19] , \AHB_IF_0_DATAOUT[20] , 
        \AHB_IF_0_DATAOUT[21] , \AHB_IF_0_DATAOUT[22] , 
        \AHB_IF_0_DATAOUT[23] , \AHB_IF_0_DATAOUT[24] , 
        \AHB_IF_0_DATAOUT[25] , \AHB_IF_0_DATAOUT[26] , 
        \AHB_IF_0_DATAOUT[27] , \AHB_IF_0_DATAOUT[28] , 
        \AHB_IF_0_DATAOUT[29] , \AHB_IF_0_DATAOUT[30] , 
        \AHB_IF_0_DATAOUT[31] , \AHB_IF_0_BIF_1_HADDR[2] , 
        \AHB_IF_0_BIF_1_HADDR[3] , \AHB_IF_0_BIF_1_HADDR[4] , 
        \AHB_IF_0_BIF_1_HADDR[5] , \AHB_IF_0_BIF_1_HADDR[6] , 
        \AHB_IF_0_BIF_1_HADDR[7] , \AHB_IF_0_BIF_1_HADDR[8] , 
        \AHB_IF_0_BIF_1_HADDR[9] , \AHB_IF_0_BIF_1_HADDR[10] , 
        \AHB_IF_0_BIF_1_HADDR[11] , \AHB_IF_0_BIF_1_HADDR[12] , 
        \AHB_IF_0_BIF_1_HADDR[13] , \AHB_IF_0_BIF_1_HADDR[14] , 
        \AHB_IF_0_BIF_1_HADDR[15] , \AHB_IF_0_BIF_1_HADDR[16] , 
        \AHB_IF_0_BIF_1_HADDR[17] , \AHB_IF_0_BIF_1_HADDR[18] , 
        \AHB_IF_0_BIF_1_HADDR[19] , \AHB_IF_0_BIF_1_HADDR[20] , 
        \AHB_IF_0_BIF_1_HADDR[21] , \AHB_IF_0_BIF_1_HADDR[22] , 
        \AHB_IF_0_BIF_1_HADDR[23] , \AHB_IF_0_BIF_1_HADDR[24] , 
        \AHB_IF_0_BIF_1_HADDR[25] , \AHB_IF_0_BIF_1_HADDR[26] , 
        \AHB_IF_0_BIF_1_HADDR[27] , \AHB_IF_0_BIF_1_HADDR[28] , 
        \AHB_IF_0_BIF_1_HADDR[29] , \AHB_IF_0_BIF_1_HADDR[30] , 
        \AHB_IF_0_BIF_1_HADDR[31] , \AHB_IF_0_BIF_1_HTRANS[1] , 
        AHB_IF_0_BIF_1_HWRITE, \AHB_IF_0_BIF_1_HWDATA[0] , 
        \AHB_IF_0_BIF_1_HWDATA[1] , \AHB_IF_0_BIF_1_HWDATA[2] , 
        \AHB_IF_0_BIF_1_HWDATA[3] , \AHB_IF_0_BIF_1_HWDATA[4] , 
        \AHB_IF_0_BIF_1_HWDATA[5] , \AHB_IF_0_BIF_1_HWDATA[6] , 
        \AHB_IF_0_BIF_1_HWDATA[7] , \AHB_IF_0_BIF_1_HWDATA[8] , 
        \AHB_IF_0_BIF_1_HWDATA[9] , \AHB_IF_0_BIF_1_HWDATA[10] , 
        \AHB_IF_0_BIF_1_HWDATA[11] , \AHB_IF_0_BIF_1_HWDATA[12] , 
        \AHB_IF_0_BIF_1_HWDATA[13] , \AHB_IF_0_BIF_1_HWDATA[14] , 
        \AHB_IF_0_BIF_1_HWDATA[15] , \AHB_IF_0_BIF_1_HWDATA[16] , 
        \AHB_IF_0_BIF_1_HWDATA[17] , \AHB_IF_0_BIF_1_HWDATA[18] , 
        \AHB_IF_0_BIF_1_HWDATA[19] , \AHB_IF_0_BIF_1_HWDATA[20] , 
        \AHB_IF_0_BIF_1_HWDATA[21] , \AHB_IF_0_BIF_1_HWDATA[22] , 
        \AHB_IF_0_BIF_1_HWDATA[23] , \AHB_IF_0_BIF_1_HWDATA[24] , 
        \AHB_IF_0_BIF_1_HWDATA[25] , \AHB_IF_0_BIF_1_HWDATA[26] , 
        \AHB_IF_0_BIF_1_HWDATA[27] , \AHB_IF_0_BIF_1_HWDATA[28] , 
        \AHB_IF_0_BIF_1_HWDATA[29] , \AHB_IF_0_BIF_1_HWDATA[30] , 
        \AHB_IF_0_BIF_1_HWDATA[31] , \AHB_IF_0_BIF_1_HRDATA[0] , 
        \AHB_IF_0_BIF_1_HRDATA[1] , \AHB_IF_0_BIF_1_HRDATA[2] , 
        \AHB_IF_0_BIF_1_HRDATA[3] , \AHB_IF_0_BIF_1_HRDATA[4] , 
        \AHB_IF_0_BIF_1_HRDATA[5] , \AHB_IF_0_BIF_1_HRDATA[6] , 
        \AHB_IF_0_BIF_1_HRDATA[7] , \AHB_IF_0_BIF_1_HRDATA[8] , 
        \AHB_IF_0_BIF_1_HRDATA[9] , \AHB_IF_0_BIF_1_HRDATA[10] , 
        \AHB_IF_0_BIF_1_HRDATA[11] , \AHB_IF_0_BIF_1_HRDATA[12] , 
        \AHB_IF_0_BIF_1_HRDATA[13] , \AHB_IF_0_BIF_1_HRDATA[14] , 
        \AHB_IF_0_BIF_1_HRDATA[15] , \AHB_IF_0_BIF_1_HRDATA[16] , 
        \AHB_IF_0_BIF_1_HRDATA[17] , \AHB_IF_0_BIF_1_HRDATA[18] , 
        \AHB_IF_0_BIF_1_HRDATA[19] , \AHB_IF_0_BIF_1_HRDATA[20] , 
        \AHB_IF_0_BIF_1_HRDATA[21] , \AHB_IF_0_BIF_1_HRDATA[22] , 
        \AHB_IF_0_BIF_1_HRDATA[23] , \AHB_IF_0_BIF_1_HRDATA[24] , 
        \AHB_IF_0_BIF_1_HRDATA[25] , \AHB_IF_0_BIF_1_HRDATA[26] , 
        \AHB_IF_0_BIF_1_HRDATA[27] , \AHB_IF_0_BIF_1_HRDATA[28] , 
        \AHB_IF_0_BIF_1_HRDATA[29] , \AHB_IF_0_BIF_1_HRDATA[30] , 
        \AHB_IF_0_BIF_1_HRDATA[31] , AHB_IF_0_AHB_BUSY, AHB_IF_0_VALID, 
        eSRAM_eNVM_RW_0_ram_wen, \eSRAM_eNVM_RW_0_ram_waddr[0] , 
        \eSRAM_eNVM_RW_0_ram_waddr[1] , \eSRAM_eNVM_RW_0_ram_waddr[2] , 
        \eSRAM_eNVM_RW_0_ram_waddr[3] , \eSRAM_eNVM_RW_0_ram_waddr[4] , 
        \eSRAM_eNVM_RW_0_ram_wdata[0] , \eSRAM_eNVM_RW_0_ram_wdata[1] , 
        \eSRAM_eNVM_RW_0_ram_wdata[2] , \eSRAM_eNVM_RW_0_ram_wdata[3] , 
        \eSRAM_eNVM_RW_0_ram_wdata[4] , \eSRAM_eNVM_RW_0_ram_wdata[5] , 
        \eSRAM_eNVM_RW_0_ram_wdata[6] , \eSRAM_eNVM_RW_0_ram_wdata[7] , 
        \eSRAM_eNVM_RW_0_ram_wdata[8] , \eSRAM_eNVM_RW_0_ram_wdata[9] , 
        \eSRAM_eNVM_RW_0_ram_wdata[10] , 
        \eSRAM_eNVM_RW_0_ram_wdata[11] , 
        \eSRAM_eNVM_RW_0_ram_wdata[12] , 
        \eSRAM_eNVM_RW_0_ram_wdata[13] , 
        \eSRAM_eNVM_RW_0_ram_wdata[14] , 
        \eSRAM_eNVM_RW_0_ram_wdata[15] , 
        \eSRAM_eNVM_RW_0_ram_wdata[16] , 
        \eSRAM_eNVM_RW_0_ram_wdata[17] , 
        \eSRAM_eNVM_RW_0_ram_wdata[18] , 
        \eSRAM_eNVM_RW_0_ram_wdata[19] , 
        \eSRAM_eNVM_RW_0_ram_wdata[20] , 
        \eSRAM_eNVM_RW_0_ram_wdata[21] , 
        \eSRAM_eNVM_RW_0_ram_wdata[22] , 
        \eSRAM_eNVM_RW_0_ram_wdata[23] , 
        \eSRAM_eNVM_RW_0_ram_wdata[24] , 
        \eSRAM_eNVM_RW_0_ram_wdata[25] , 
        \eSRAM_eNVM_RW_0_ram_wdata[26] , 
        \eSRAM_eNVM_RW_0_ram_wdata[27] , 
        \eSRAM_eNVM_RW_0_ram_wdata[28] , 
        \eSRAM_eNVM_RW_0_ram_wdata[29] , 
        \eSRAM_eNVM_RW_0_ram_wdata[30] , 
        \eSRAM_eNVM_RW_0_ram_wdata[31] , CLKOUT_1, MOSI_1, 
        \SPI_Master_0.state[0] , 
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState , 
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMNextState , 
        FAB_RESET_N_c, MISO_c, PWRITE_c, start_esram_c, CS_c, 
        \PRDATA_c[0] , \PRDATA_c[1] , \PRDATA_c[2] , \PRDATA_c[3] , 
        \PRDATA_c[4] , \PRDATA_c[5] , \PRDATA_c[6] , \PRDATA_c[7] , 
        \PRDATA_c[8] , \PRDATA_c[9] , \PRDATA_c[10] , \PRDATA_c[11] , 
        \PRDATA_c[12] , \PRDATA_c[13] , \PRDATA_c[14] , \PRDATA_c[15] , 
        \PRDATA_c[16] , \PRDATA_c[17] , \PRDATA_c[18] , \PRDATA_c[19] , 
        \PRDATA_c[20] , \PRDATA_c[21] , \PRDATA_c[22] , \PRDATA_c[23] , 
        \PRDATA_c[24] , \PRDATA_c[25] , \PRDATA_c[26] , \PRDATA_c[27] , 
        \PRDATA_c[28] , \PRDATA_c[29] , \PRDATA_c[30] , \PRDATA_c[31] , 
        \RD_c[0] , \RD_c[1] , \RD_c[2] , \RD_c[3] , \RD_c[4] , 
        \RD_c[5] , \RD_c[6] , \RD_c[7] , ss_n_c, N_546, N_53, 
        \eSRAM_eNVM_RW_0_ADDR[3] , \eSRAM_eNVM_RW_0_ADDR[4] , 
        \eSRAM_eNVM_RW_0_ADDR[5] , \eSRAM_eNVM_RW_0_ADDR[6] , 
        \eSRAM_eNVM_RW_0_ADDR[7] , \eSRAM_eNVM_RW_0_ADDR[8] , 
        \eSRAM_eNVM_RW_0_ADDR[9] , \eSRAM_eNVM_RW_0_ADDR[10] , 
        \eSRAM_eNVM_RW_0_ADDR[11] , \eSRAM_eNVM_RW_0_ADDR[12] , 
        \eSRAM_eNVM_RW_0_ADDR[13] , \eSRAM_eNVM_RW_0_ADDR[14] , 
        \eSRAM_eNVM_RW_0_ADDR[15] , \eSRAM_eNVM_RW_0_ADDR[16] , 
        \eSRAM_eNVM_RW_0_ADDR[17] , \eSRAM_eNVM_RW_0_ADDR[18] , 
        \eSRAM_eNVM_RW_0_ADDR[19] , \eSRAM_eNVM_RW_0_ADDR[20] , 
        \eSRAM_eNVM_RW_0_ADDR[21] , \eSRAM_eNVM_RW_0_ADDR[22] , 
        \eSRAM_eNVM_RW_0_ADDR[23] , \eSRAM_eNVM_RW_0_ADDR[24] , 
        \eSRAM_eNVM_RW_0_ADDR[25] , \eSRAM_eNVM_RW_0_ADDR[26] , 
        \eSRAM_eNVM_RW_0_ADDR[27] , \eSRAM_eNVM_RW_0_ADDR[28] , 
        \eSRAM_eNVM_RW_0_ADDR[29] , \eSRAM_eNVM_RW_0_ADDR[30] , 
        \eSRAM_eNVM_RW_0_ADDR[31] , \eSRAM_eNVM_RW_0_DATAOUT[1] , 
        \eSRAM_eNVM_RW_0_DATAOUT[2] , \eSRAM_eNVM_RW_0_DATAOUT[3] , 
        \eSRAM_eNVM_RW_0_DATAOUT[4] , \eSRAM_eNVM_RW_0_DATAOUT[5] , 
        \eSRAM_eNVM_RW_0_DATAOUT[6] , \eSRAM_eNVM_RW_0_DATAOUT[7] , 
        \eSRAM_eNVM_RW_0_DATAOUT[8] , \eSRAM_eNVM_RW_0_DATAOUT[9] , 
        \eSRAM_eNVM_RW_0_DATAOUT[10] , \eSRAM_eNVM_RW_0_DATAOUT[11] , 
        \eSRAM_eNVM_RW_0_DATAOUT[12] , \eSRAM_eNVM_RW_0_DATAOUT[13] , 
        \eSRAM_eNVM_RW_0_DATAOUT[14] , \eSRAM_eNVM_RW_0_DATAOUT[15] , 
        \eSRAM_eNVM_RW_0_DATAOUT[16] , \eSRAM_eNVM_RW_0_DATAOUT[17] , 
        \eSRAM_eNVM_RW_0_DATAOUT[18] , \eSRAM_eNVM_RW_0_DATAOUT[19] , 
        \eSRAM_eNVM_RW_0_DATAOUT[20] , \eSRAM_eNVM_RW_0_DATAOUT[21] , 
        \eSRAM_eNVM_RW_0_DATAOUT[22] , \eSRAM_eNVM_RW_0_DATAOUT[23] , 
        \eSRAM_eNVM_RW_0_DATAOUT[24] , \eSRAM_eNVM_RW_0_DATAOUT[25] , 
        \eSRAM_eNVM_RW_0_DATAOUT[26] , \eSRAM_eNVM_RW_0_DATAOUT[27] , 
        \eSRAM_eNVM_RW_0_DATAOUT[28] , \eSRAM_eNVM_RW_0_DATAOUT[29] , 
        \eSRAM_eNVM_RW_0_DATAOUT[30] , \eSRAM_eNVM_RW_0_DATAOUT[31] , 
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.HREADY_M_0_iv_i_0 , 
        MOSI_cl, CLKOUT_cl;
    
    eSRAM_eNVM_access_top_TPSRAM_0_TPSRAM TPSRAM_0 (.RD_c({\RD_c[7] , 
        \RD_c[6] , \RD_c[5] , \RD_c[4] , \RD_c[3] , \RD_c[2] , 
        \RD_c[1] , \RD_c[0] }), .eSRAM_eNVM_RW_0_ram_wdata({
        \eSRAM_eNVM_RW_0_ram_wdata[31] , 
        \eSRAM_eNVM_RW_0_ram_wdata[30] , 
        \eSRAM_eNVM_RW_0_ram_wdata[29] , 
        \eSRAM_eNVM_RW_0_ram_wdata[28] , 
        \eSRAM_eNVM_RW_0_ram_wdata[27] , 
        \eSRAM_eNVM_RW_0_ram_wdata[26] , 
        \eSRAM_eNVM_RW_0_ram_wdata[25] , 
        \eSRAM_eNVM_RW_0_ram_wdata[24] , 
        \eSRAM_eNVM_RW_0_ram_wdata[23] , 
        \eSRAM_eNVM_RW_0_ram_wdata[22] , 
        \eSRAM_eNVM_RW_0_ram_wdata[21] , 
        \eSRAM_eNVM_RW_0_ram_wdata[20] , 
        \eSRAM_eNVM_RW_0_ram_wdata[19] , 
        \eSRAM_eNVM_RW_0_ram_wdata[18] , 
        \eSRAM_eNVM_RW_0_ram_wdata[17] , 
        \eSRAM_eNVM_RW_0_ram_wdata[16] , 
        \eSRAM_eNVM_RW_0_ram_wdata[15] , 
        \eSRAM_eNVM_RW_0_ram_wdata[14] , 
        \eSRAM_eNVM_RW_0_ram_wdata[13] , 
        \eSRAM_eNVM_RW_0_ram_wdata[12] , 
        \eSRAM_eNVM_RW_0_ram_wdata[11] , 
        \eSRAM_eNVM_RW_0_ram_wdata[10] , 
        \eSRAM_eNVM_RW_0_ram_wdata[9] , \eSRAM_eNVM_RW_0_ram_wdata[8] , 
        \eSRAM_eNVM_RW_0_ram_wdata[7] , \eSRAM_eNVM_RW_0_ram_wdata[6] , 
        \eSRAM_eNVM_RW_0_ram_wdata[5] , \eSRAM_eNVM_RW_0_ram_wdata[4] , 
        \eSRAM_eNVM_RW_0_ram_wdata[3] , \eSRAM_eNVM_RW_0_ram_wdata[2] , 
        \eSRAM_eNVM_RW_0_ram_wdata[1] , \eSRAM_eNVM_RW_0_ram_wdata[0] })
        , .eSRAM_eNVM_RW_0_ram_waddr({\eSRAM_eNVM_RW_0_ram_waddr[4] , 
        \eSRAM_eNVM_RW_0_ram_waddr[3] , \eSRAM_eNVM_RW_0_ram_waddr[2] , 
        \eSRAM_eNVM_RW_0_ram_waddr[1] , \eSRAM_eNVM_RW_0_ram_waddr[0] })
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .eSRAM_eNVM_RW_0_ram_wen(eSRAM_eNVM_RW_0_ram_wen));
    eSRAM_eNVM_access eSRAM_eNVM_access_0 (.AHB_IF_0_BIF_1_HADDR({
        \AHB_IF_0_BIF_1_HADDR[31] , \AHB_IF_0_BIF_1_HADDR[30] , 
        \AHB_IF_0_BIF_1_HADDR[29] , \AHB_IF_0_BIF_1_HADDR[28] , 
        \AHB_IF_0_BIF_1_HADDR[27] , \AHB_IF_0_BIF_1_HADDR[26] , 
        \AHB_IF_0_BIF_1_HADDR[25] , \AHB_IF_0_BIF_1_HADDR[24] , 
        \AHB_IF_0_BIF_1_HADDR[23] , \AHB_IF_0_BIF_1_HADDR[22] , 
        \AHB_IF_0_BIF_1_HADDR[21] , \AHB_IF_0_BIF_1_HADDR[20] , 
        \AHB_IF_0_BIF_1_HADDR[19] , \AHB_IF_0_BIF_1_HADDR[18] , 
        \AHB_IF_0_BIF_1_HADDR[17] , \AHB_IF_0_BIF_1_HADDR[16] , 
        \AHB_IF_0_BIF_1_HADDR[15] , \AHB_IF_0_BIF_1_HADDR[14] , 
        \AHB_IF_0_BIF_1_HADDR[13] , \AHB_IF_0_BIF_1_HADDR[12] , 
        \AHB_IF_0_BIF_1_HADDR[11] , \AHB_IF_0_BIF_1_HADDR[10] , 
        \AHB_IF_0_BIF_1_HADDR[9] , \AHB_IF_0_BIF_1_HADDR[8] , 
        \AHB_IF_0_BIF_1_HADDR[7] , \AHB_IF_0_BIF_1_HADDR[6] , 
        \AHB_IF_0_BIF_1_HADDR[5] , \AHB_IF_0_BIF_1_HADDR[4] , 
        \AHB_IF_0_BIF_1_HADDR[3] , \AHB_IF_0_BIF_1_HADDR[2] }), 
        .AHB_IF_0_BIF_1_HTRANS({\AHB_IF_0_BIF_1_HTRANS[1] }), 
        .AHB_IF_0_BIF_1_HWDATA({\AHB_IF_0_BIF_1_HWDATA[31] , 
        \AHB_IF_0_BIF_1_HWDATA[30] , \AHB_IF_0_BIF_1_HWDATA[29] , 
        \AHB_IF_0_BIF_1_HWDATA[28] , \AHB_IF_0_BIF_1_HWDATA[27] , 
        \AHB_IF_0_BIF_1_HWDATA[26] , \AHB_IF_0_BIF_1_HWDATA[25] , 
        \AHB_IF_0_BIF_1_HWDATA[24] , \AHB_IF_0_BIF_1_HWDATA[23] , 
        \AHB_IF_0_BIF_1_HWDATA[22] , \AHB_IF_0_BIF_1_HWDATA[21] , 
        \AHB_IF_0_BIF_1_HWDATA[20] , \AHB_IF_0_BIF_1_HWDATA[19] , 
        \AHB_IF_0_BIF_1_HWDATA[18] , \AHB_IF_0_BIF_1_HWDATA[17] , 
        \AHB_IF_0_BIF_1_HWDATA[16] , \AHB_IF_0_BIF_1_HWDATA[15] , 
        \AHB_IF_0_BIF_1_HWDATA[14] , \AHB_IF_0_BIF_1_HWDATA[13] , 
        \AHB_IF_0_BIF_1_HWDATA[12] , \AHB_IF_0_BIF_1_HWDATA[11] , 
        \AHB_IF_0_BIF_1_HWDATA[10] , \AHB_IF_0_BIF_1_HWDATA[9] , 
        \AHB_IF_0_BIF_1_HWDATA[8] , \AHB_IF_0_BIF_1_HWDATA[7] , 
        \AHB_IF_0_BIF_1_HWDATA[6] , \AHB_IF_0_BIF_1_HWDATA[5] , 
        \AHB_IF_0_BIF_1_HWDATA[4] , \AHB_IF_0_BIF_1_HWDATA[3] , 
        \AHB_IF_0_BIF_1_HWDATA[2] , \AHB_IF_0_BIF_1_HWDATA[1] , 
        \AHB_IF_0_BIF_1_HWDATA[0] }), .AHB_IF_0_BIF_1_HRDATA({
        \AHB_IF_0_BIF_1_HRDATA[31] , \AHB_IF_0_BIF_1_HRDATA[30] , 
        \AHB_IF_0_BIF_1_HRDATA[29] , \AHB_IF_0_BIF_1_HRDATA[28] , 
        \AHB_IF_0_BIF_1_HRDATA[27] , \AHB_IF_0_BIF_1_HRDATA[26] , 
        \AHB_IF_0_BIF_1_HRDATA[25] , \AHB_IF_0_BIF_1_HRDATA[24] , 
        \AHB_IF_0_BIF_1_HRDATA[23] , \AHB_IF_0_BIF_1_HRDATA[22] , 
        \AHB_IF_0_BIF_1_HRDATA[21] , \AHB_IF_0_BIF_1_HRDATA[20] , 
        \AHB_IF_0_BIF_1_HRDATA[19] , \AHB_IF_0_BIF_1_HRDATA[18] , 
        \AHB_IF_0_BIF_1_HRDATA[17] , \AHB_IF_0_BIF_1_HRDATA[16] , 
        \AHB_IF_0_BIF_1_HRDATA[15] , \AHB_IF_0_BIF_1_HRDATA[14] , 
        \AHB_IF_0_BIF_1_HRDATA[13] , \AHB_IF_0_BIF_1_HRDATA[12] , 
        \AHB_IF_0_BIF_1_HRDATA[11] , \AHB_IF_0_BIF_1_HRDATA[10] , 
        \AHB_IF_0_BIF_1_HRDATA[9] , \AHB_IF_0_BIF_1_HRDATA[8] , 
        \AHB_IF_0_BIF_1_HRDATA[7] , \AHB_IF_0_BIF_1_HRDATA[6] , 
        \AHB_IF_0_BIF_1_HRDATA[5] , \AHB_IF_0_BIF_1_HRDATA[4] , 
        \AHB_IF_0_BIF_1_HRDATA[3] , \AHB_IF_0_BIF_1_HRDATA[2] , 
        \AHB_IF_0_BIF_1_HRDATA[1] , \AHB_IF_0_BIF_1_HRDATA[0] }), 
        .DEVRST_N(DEVRST_N), .eSRAM_eNVM_access_0_FIC_0_CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .AHB_IF_0_BIF_1_HWRITE(AHB_IF_0_BIF_1_HWRITE), 
        .defSlaveSMCurrentState(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState )
        , .defSlaveSMNextState(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMNextState )
        , .N_53(N_53), .N_546(N_546), .HREADY_M_0_iv_i_0(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.HREADY_M_0_iv_i_0 )
        , .FAB_RESET_N_c(FAB_RESET_N_c));
    OUTBUF \PRDATA_obuf[14]  (.D(\PRDATA_c[14] ), .PAD(PRDATA[14]));
    OUTBUF \PRDATA_obuf[27]  (.D(\PRDATA_c[27] ), .PAD(PRDATA[27]));
    INBUF start_esram_ibuf (.PAD(start_esram), .Y(start_esram_c));
    OUTBUF \PRDATA_obuf[18]  (.D(\PRDATA_c[18] ), .PAD(PRDATA[18]));
    OUTBUF \PRDATA_obuf[29]  (.D(\PRDATA_c[29] ), .PAD(PRDATA[29]));
    OUTBUF \RD_obuf[2]  (.D(\RD_c[2] ), .PAD(RD[2]));
    OUTBUF \RD_obuf[6]  (.D(\RD_c[6] ), .PAD(RD[6]));
    OUTBUF \PRDATA_obuf[8]  (.D(\PRDATA_c[8] ), .PAD(PRDATA[8]));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF \PRDATA_obuf[20]  (.D(\PRDATA_c[20] ), .PAD(PRDATA[20]));
    OUTBUF \PRDATA_obuf[11]  (.D(\PRDATA_c[11] ), .PAD(PRDATA[11]));
    INBUF MISO_ibuf (.PAD(MISO), .Y(MISO_c));
    OUTBUF ss_n_obuf (.D(ss_n_c), .PAD(ss_n));
    OUTBUF \PRDATA_obuf[22]  (.D(\PRDATA_c[22] ), .PAD(PRDATA[22]));
    OUTBUF \RD_obuf[3]  (.D(\RD_c[3] ), .PAD(RD[3]));
    eSRAM_eNVM_RW eSRAM_eNVM_RW_0 (.eSRAM_eNVM_RW_0_ram_waddr({
        \eSRAM_eNVM_RW_0_ram_waddr[4] , \eSRAM_eNVM_RW_0_ram_waddr[3] , 
        \eSRAM_eNVM_RW_0_ram_waddr[2] , \eSRAM_eNVM_RW_0_ram_waddr[1] , 
        \eSRAM_eNVM_RW_0_ram_waddr[0] }), .eSRAM_eNVM_RW_0_ram_wdata({
        \eSRAM_eNVM_RW_0_ram_wdata[31] , 
        \eSRAM_eNVM_RW_0_ram_wdata[30] , 
        \eSRAM_eNVM_RW_0_ram_wdata[29] , 
        \eSRAM_eNVM_RW_0_ram_wdata[28] , 
        \eSRAM_eNVM_RW_0_ram_wdata[27] , 
        \eSRAM_eNVM_RW_0_ram_wdata[26] , 
        \eSRAM_eNVM_RW_0_ram_wdata[25] , 
        \eSRAM_eNVM_RW_0_ram_wdata[24] , 
        \eSRAM_eNVM_RW_0_ram_wdata[23] , 
        \eSRAM_eNVM_RW_0_ram_wdata[22] , 
        \eSRAM_eNVM_RW_0_ram_wdata[21] , 
        \eSRAM_eNVM_RW_0_ram_wdata[20] , 
        \eSRAM_eNVM_RW_0_ram_wdata[19] , 
        \eSRAM_eNVM_RW_0_ram_wdata[18] , 
        \eSRAM_eNVM_RW_0_ram_wdata[17] , 
        \eSRAM_eNVM_RW_0_ram_wdata[16] , 
        \eSRAM_eNVM_RW_0_ram_wdata[15] , 
        \eSRAM_eNVM_RW_0_ram_wdata[14] , 
        \eSRAM_eNVM_RW_0_ram_wdata[13] , 
        \eSRAM_eNVM_RW_0_ram_wdata[12] , 
        \eSRAM_eNVM_RW_0_ram_wdata[11] , 
        \eSRAM_eNVM_RW_0_ram_wdata[10] , 
        \eSRAM_eNVM_RW_0_ram_wdata[9] , \eSRAM_eNVM_RW_0_ram_wdata[8] , 
        \eSRAM_eNVM_RW_0_ram_wdata[7] , \eSRAM_eNVM_RW_0_ram_wdata[6] , 
        \eSRAM_eNVM_RW_0_ram_wdata[5] , \eSRAM_eNVM_RW_0_ram_wdata[4] , 
        \eSRAM_eNVM_RW_0_ram_wdata[3] , \eSRAM_eNVM_RW_0_ram_wdata[2] , 
        \eSRAM_eNVM_RW_0_ram_wdata[1] , \eSRAM_eNVM_RW_0_ram_wdata[0] })
        , .AHB_IF_0_DATAOUT({\AHB_IF_0_DATAOUT[31] , 
        \AHB_IF_0_DATAOUT[30] , \AHB_IF_0_DATAOUT[29] , 
        \AHB_IF_0_DATAOUT[28] , \AHB_IF_0_DATAOUT[27] , 
        \AHB_IF_0_DATAOUT[26] , \AHB_IF_0_DATAOUT[25] , 
        \AHB_IF_0_DATAOUT[24] , \AHB_IF_0_DATAOUT[23] , 
        \AHB_IF_0_DATAOUT[22] , \AHB_IF_0_DATAOUT[21] , 
        \AHB_IF_0_DATAOUT[20] , \AHB_IF_0_DATAOUT[19] , 
        \AHB_IF_0_DATAOUT[18] , \AHB_IF_0_DATAOUT[17] , 
        \AHB_IF_0_DATAOUT[16] , \AHB_IF_0_DATAOUT[15] , 
        \AHB_IF_0_DATAOUT[14] , \AHB_IF_0_DATAOUT[13] , 
        \AHB_IF_0_DATAOUT[12] , \AHB_IF_0_DATAOUT[11] , 
        \AHB_IF_0_DATAOUT[10] , \AHB_IF_0_DATAOUT[9] , 
        \AHB_IF_0_DATAOUT[8] , \AHB_IF_0_DATAOUT[7] , 
        \AHB_IF_0_DATAOUT[6] , \AHB_IF_0_DATAOUT[5] , 
        \AHB_IF_0_DATAOUT[4] , \AHB_IF_0_DATAOUT[3] , 
        \AHB_IF_0_DATAOUT[2] , \AHB_IF_0_DATAOUT[1] , 
        \AHB_IF_0_DATAOUT[0] }), .state({\SPI_Master_0.state[0] }), 
        .eSRAM_eNVM_RW_0_ADDR({\eSRAM_eNVM_RW_0_ADDR[31] , 
        \eSRAM_eNVM_RW_0_ADDR[30] , \eSRAM_eNVM_RW_0_ADDR[29] , 
        \eSRAM_eNVM_RW_0_ADDR[28] , \eSRAM_eNVM_RW_0_ADDR[27] , 
        \eSRAM_eNVM_RW_0_ADDR[26] , \eSRAM_eNVM_RW_0_ADDR[25] , 
        \eSRAM_eNVM_RW_0_ADDR[24] , \eSRAM_eNVM_RW_0_ADDR[23] , 
        \eSRAM_eNVM_RW_0_ADDR[22] , \eSRAM_eNVM_RW_0_ADDR[21] , 
        \eSRAM_eNVM_RW_0_ADDR[20] , \eSRAM_eNVM_RW_0_ADDR[19] , 
        \eSRAM_eNVM_RW_0_ADDR[18] , \eSRAM_eNVM_RW_0_ADDR[17] , 
        \eSRAM_eNVM_RW_0_ADDR[16] , \eSRAM_eNVM_RW_0_ADDR[15] , 
        \eSRAM_eNVM_RW_0_ADDR[14] , \eSRAM_eNVM_RW_0_ADDR[13] , 
        \eSRAM_eNVM_RW_0_ADDR[12] , \eSRAM_eNVM_RW_0_ADDR[11] , 
        \eSRAM_eNVM_RW_0_ADDR[10] , \eSRAM_eNVM_RW_0_ADDR[9] , 
        \eSRAM_eNVM_RW_0_ADDR[8] , \eSRAM_eNVM_RW_0_ADDR[7] , 
        \eSRAM_eNVM_RW_0_ADDR[6] , \eSRAM_eNVM_RW_0_ADDR[5] , 
        \eSRAM_eNVM_RW_0_ADDR[4] , \eSRAM_eNVM_RW_0_ADDR[3] , 
        \eSRAM_eNVM_RW_0_ADDR[2] }), .eSRAM_eNVM_RW_0_DATAOUT({
        \eSRAM_eNVM_RW_0_DATAOUT[31] , \eSRAM_eNVM_RW_0_DATAOUT[30] , 
        \eSRAM_eNVM_RW_0_DATAOUT[29] , \eSRAM_eNVM_RW_0_DATAOUT[28] , 
        \eSRAM_eNVM_RW_0_DATAOUT[27] , \eSRAM_eNVM_RW_0_DATAOUT[26] , 
        \eSRAM_eNVM_RW_0_DATAOUT[25] , \eSRAM_eNVM_RW_0_DATAOUT[24] , 
        \eSRAM_eNVM_RW_0_DATAOUT[23] , \eSRAM_eNVM_RW_0_DATAOUT[22] , 
        \eSRAM_eNVM_RW_0_DATAOUT[21] , \eSRAM_eNVM_RW_0_DATAOUT[20] , 
        \eSRAM_eNVM_RW_0_DATAOUT[19] , \eSRAM_eNVM_RW_0_DATAOUT[18] , 
        \eSRAM_eNVM_RW_0_DATAOUT[17] , \eSRAM_eNVM_RW_0_DATAOUT[16] , 
        \eSRAM_eNVM_RW_0_DATAOUT[15] , \eSRAM_eNVM_RW_0_DATAOUT[14] , 
        \eSRAM_eNVM_RW_0_DATAOUT[13] , \eSRAM_eNVM_RW_0_DATAOUT[12] , 
        \eSRAM_eNVM_RW_0_DATAOUT[11] , \eSRAM_eNVM_RW_0_DATAOUT[10] , 
        \eSRAM_eNVM_RW_0_DATAOUT[9] , \eSRAM_eNVM_RW_0_DATAOUT[8] , 
        \eSRAM_eNVM_RW_0_DATAOUT[7] , \eSRAM_eNVM_RW_0_DATAOUT[6] , 
        \eSRAM_eNVM_RW_0_DATAOUT[5] , \eSRAM_eNVM_RW_0_DATAOUT[4] , 
        \eSRAM_eNVM_RW_0_DATAOUT[3] , \eSRAM_eNVM_RW_0_DATAOUT[2] , 
        \eSRAM_eNVM_RW_0_DATAOUT[1] , \eSRAM_eNVM_RW_0_DATAOUT[0] }), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .eSRAM_eNVM_access_0_FIC_0_CLK(eSRAM_eNVM_access_0_FIC_0_CLK)
        , .eSRAM_eNVM_RW_0_WRITE(eSRAM_eNVM_RW_0_WRITE), 
        .eSRAM_eNVM_RW_0_READ(eSRAM_eNVM_RW_0_READ), 
        .eSRAM_eNVM_RW_0_ram_wen(eSRAM_eNVM_RW_0_ram_wen), 
        .start_esram_c(start_esram_c), .AHB_IF_0_AHB_BUSY(
        AHB_IF_0_AHB_BUSY), .AHB_IF_0_VALID(AHB_IF_0_VALID));
    OUTBUF \PRDATA_obuf[31]  (.D(\PRDATA_c[31] ), .PAD(PRDATA[31]));
    OUTBUF \PRDATA_obuf[26]  (.D(\PRDATA_c[26] ), .PAD(PRDATA[26]));
    OUTBUF \PRDATA_obuf[25]  (.D(\PRDATA_c[25] ), .PAD(PRDATA[25]));
    OUTBUF \PRDATA_obuf[1]  (.D(\PRDATA_c[1] ), .PAD(PRDATA[1]));
    TRIBUFF MOSI_obuft (.D(MOSI_1), .E(MOSI_cl), .PAD(MOSI));
    AHB_IF_0s_1s_2s_3s_4294967292s_4294967293s_4294967294s_0s_1_layer0 
        AHB_IF_0 (.eSRAM_eNVM_RW_0_DATAOUT({
        \eSRAM_eNVM_RW_0_DATAOUT[31] , \eSRAM_eNVM_RW_0_DATAOUT[30] , 
        \eSRAM_eNVM_RW_0_DATAOUT[29] , \eSRAM_eNVM_RW_0_DATAOUT[28] , 
        \eSRAM_eNVM_RW_0_DATAOUT[27] , \eSRAM_eNVM_RW_0_DATAOUT[26] , 
        \eSRAM_eNVM_RW_0_DATAOUT[25] , \eSRAM_eNVM_RW_0_DATAOUT[24] , 
        \eSRAM_eNVM_RW_0_DATAOUT[23] , \eSRAM_eNVM_RW_0_DATAOUT[22] , 
        \eSRAM_eNVM_RW_0_DATAOUT[21] , \eSRAM_eNVM_RW_0_DATAOUT[20] , 
        \eSRAM_eNVM_RW_0_DATAOUT[19] , \eSRAM_eNVM_RW_0_DATAOUT[18] , 
        \eSRAM_eNVM_RW_0_DATAOUT[17] , \eSRAM_eNVM_RW_0_DATAOUT[16] , 
        \eSRAM_eNVM_RW_0_DATAOUT[15] , \eSRAM_eNVM_RW_0_DATAOUT[14] , 
        \eSRAM_eNVM_RW_0_DATAOUT[13] , \eSRAM_eNVM_RW_0_DATAOUT[12] , 
        \eSRAM_eNVM_RW_0_DATAOUT[11] , \eSRAM_eNVM_RW_0_DATAOUT[10] , 
        \eSRAM_eNVM_RW_0_DATAOUT[9] , \eSRAM_eNVM_RW_0_DATAOUT[8] , 
        \eSRAM_eNVM_RW_0_DATAOUT[7] , \eSRAM_eNVM_RW_0_DATAOUT[6] , 
        \eSRAM_eNVM_RW_0_DATAOUT[5] , \eSRAM_eNVM_RW_0_DATAOUT[4] , 
        \eSRAM_eNVM_RW_0_DATAOUT[3] , \eSRAM_eNVM_RW_0_DATAOUT[2] , 
        \eSRAM_eNVM_RW_0_DATAOUT[1] , \eSRAM_eNVM_RW_0_DATAOUT[0] }), 
        .AHB_IF_0_DATAOUT({\AHB_IF_0_DATAOUT[31] , 
        \AHB_IF_0_DATAOUT[30] , \AHB_IF_0_DATAOUT[29] , 
        \AHB_IF_0_DATAOUT[28] , \AHB_IF_0_DATAOUT[27] , 
        \AHB_IF_0_DATAOUT[26] , \AHB_IF_0_DATAOUT[25] , 
        \AHB_IF_0_DATAOUT[24] , \AHB_IF_0_DATAOUT[23] , 
        \AHB_IF_0_DATAOUT[22] , \AHB_IF_0_DATAOUT[21] , 
        \AHB_IF_0_DATAOUT[20] , \AHB_IF_0_DATAOUT[19] , 
        \AHB_IF_0_DATAOUT[18] , \AHB_IF_0_DATAOUT[17] , 
        \AHB_IF_0_DATAOUT[16] , \AHB_IF_0_DATAOUT[15] , 
        \AHB_IF_0_DATAOUT[14] , \AHB_IF_0_DATAOUT[13] , 
        \AHB_IF_0_DATAOUT[12] , \AHB_IF_0_DATAOUT[11] , 
        \AHB_IF_0_DATAOUT[10] , \AHB_IF_0_DATAOUT[9] , 
        \AHB_IF_0_DATAOUT[8] , \AHB_IF_0_DATAOUT[7] , 
        \AHB_IF_0_DATAOUT[6] , \AHB_IF_0_DATAOUT[5] , 
        \AHB_IF_0_DATAOUT[4] , \AHB_IF_0_DATAOUT[3] , 
        \AHB_IF_0_DATAOUT[2] , \AHB_IF_0_DATAOUT[1] , 
        \AHB_IF_0_DATAOUT[0] }), .AHB_IF_0_BIF_1_HRDATA({
        \AHB_IF_0_BIF_1_HRDATA[31] , \AHB_IF_0_BIF_1_HRDATA[30] , 
        \AHB_IF_0_BIF_1_HRDATA[29] , \AHB_IF_0_BIF_1_HRDATA[28] , 
        \AHB_IF_0_BIF_1_HRDATA[27] , \AHB_IF_0_BIF_1_HRDATA[26] , 
        \AHB_IF_0_BIF_1_HRDATA[25] , \AHB_IF_0_BIF_1_HRDATA[24] , 
        \AHB_IF_0_BIF_1_HRDATA[23] , \AHB_IF_0_BIF_1_HRDATA[22] , 
        \AHB_IF_0_BIF_1_HRDATA[21] , \AHB_IF_0_BIF_1_HRDATA[20] , 
        \AHB_IF_0_BIF_1_HRDATA[19] , \AHB_IF_0_BIF_1_HRDATA[18] , 
        \AHB_IF_0_BIF_1_HRDATA[17] , \AHB_IF_0_BIF_1_HRDATA[16] , 
        \AHB_IF_0_BIF_1_HRDATA[15] , \AHB_IF_0_BIF_1_HRDATA[14] , 
        \AHB_IF_0_BIF_1_HRDATA[13] , \AHB_IF_0_BIF_1_HRDATA[12] , 
        \AHB_IF_0_BIF_1_HRDATA[11] , \AHB_IF_0_BIF_1_HRDATA[10] , 
        \AHB_IF_0_BIF_1_HRDATA[9] , \AHB_IF_0_BIF_1_HRDATA[8] , 
        \AHB_IF_0_BIF_1_HRDATA[7] , \AHB_IF_0_BIF_1_HRDATA[6] , 
        \AHB_IF_0_BIF_1_HRDATA[5] , \AHB_IF_0_BIF_1_HRDATA[4] , 
        \AHB_IF_0_BIF_1_HRDATA[3] , \AHB_IF_0_BIF_1_HRDATA[2] , 
        \AHB_IF_0_BIF_1_HRDATA[1] , \AHB_IF_0_BIF_1_HRDATA[0] }), 
        .AHB_IF_0_BIF_1_HWDATA({\AHB_IF_0_BIF_1_HWDATA[31] , 
        \AHB_IF_0_BIF_1_HWDATA[30] , \AHB_IF_0_BIF_1_HWDATA[29] , 
        \AHB_IF_0_BIF_1_HWDATA[28] , \AHB_IF_0_BIF_1_HWDATA[27] , 
        \AHB_IF_0_BIF_1_HWDATA[26] , \AHB_IF_0_BIF_1_HWDATA[25] , 
        \AHB_IF_0_BIF_1_HWDATA[24] , \AHB_IF_0_BIF_1_HWDATA[23] , 
        \AHB_IF_0_BIF_1_HWDATA[22] , \AHB_IF_0_BIF_1_HWDATA[21] , 
        \AHB_IF_0_BIF_1_HWDATA[20] , \AHB_IF_0_BIF_1_HWDATA[19] , 
        \AHB_IF_0_BIF_1_HWDATA[18] , \AHB_IF_0_BIF_1_HWDATA[17] , 
        \AHB_IF_0_BIF_1_HWDATA[16] , \AHB_IF_0_BIF_1_HWDATA[15] , 
        \AHB_IF_0_BIF_1_HWDATA[14] , \AHB_IF_0_BIF_1_HWDATA[13] , 
        \AHB_IF_0_BIF_1_HWDATA[12] , \AHB_IF_0_BIF_1_HWDATA[11] , 
        \AHB_IF_0_BIF_1_HWDATA[10] , \AHB_IF_0_BIF_1_HWDATA[9] , 
        \AHB_IF_0_BIF_1_HWDATA[8] , \AHB_IF_0_BIF_1_HWDATA[7] , 
        \AHB_IF_0_BIF_1_HWDATA[6] , \AHB_IF_0_BIF_1_HWDATA[5] , 
        \AHB_IF_0_BIF_1_HWDATA[4] , \AHB_IF_0_BIF_1_HWDATA[3] , 
        \AHB_IF_0_BIF_1_HWDATA[2] , \AHB_IF_0_BIF_1_HWDATA[1] , 
        \AHB_IF_0_BIF_1_HWDATA[0] }), .AHB_IF_0_BIF_1_HADDR({
        \AHB_IF_0_BIF_1_HADDR[31] , \AHB_IF_0_BIF_1_HADDR[30] , 
        \AHB_IF_0_BIF_1_HADDR[29] , \AHB_IF_0_BIF_1_HADDR[28] , 
        \AHB_IF_0_BIF_1_HADDR[27] , \AHB_IF_0_BIF_1_HADDR[26] , 
        \AHB_IF_0_BIF_1_HADDR[25] , \AHB_IF_0_BIF_1_HADDR[24] , 
        \AHB_IF_0_BIF_1_HADDR[23] , \AHB_IF_0_BIF_1_HADDR[22] , 
        \AHB_IF_0_BIF_1_HADDR[21] , \AHB_IF_0_BIF_1_HADDR[20] , 
        \AHB_IF_0_BIF_1_HADDR[19] , \AHB_IF_0_BIF_1_HADDR[18] , 
        \AHB_IF_0_BIF_1_HADDR[17] , \AHB_IF_0_BIF_1_HADDR[16] , 
        \AHB_IF_0_BIF_1_HADDR[15] , \AHB_IF_0_BIF_1_HADDR[14] , 
        \AHB_IF_0_BIF_1_HADDR[13] , \AHB_IF_0_BIF_1_HADDR[12] , 
        \AHB_IF_0_BIF_1_HADDR[11] , \AHB_IF_0_BIF_1_HADDR[10] , 
        \AHB_IF_0_BIF_1_HADDR[9] , \AHB_IF_0_BIF_1_HADDR[8] , 
        \AHB_IF_0_BIF_1_HADDR[7] , \AHB_IF_0_BIF_1_HADDR[6] , 
        \AHB_IF_0_BIF_1_HADDR[5] , \AHB_IF_0_BIF_1_HADDR[4] , 
        \AHB_IF_0_BIF_1_HADDR[3] , \AHB_IF_0_BIF_1_HADDR[2] }), 
        .AHB_IF_0_BIF_1_HTRANS({\AHB_IF_0_BIF_1_HTRANS[1] }), 
        .eSRAM_eNVM_RW_0_ADDR({\eSRAM_eNVM_RW_0_ADDR[31] , 
        \eSRAM_eNVM_RW_0_ADDR[30] , \eSRAM_eNVM_RW_0_ADDR[29] , 
        \eSRAM_eNVM_RW_0_ADDR[28] , \eSRAM_eNVM_RW_0_ADDR[27] , 
        \eSRAM_eNVM_RW_0_ADDR[26] , \eSRAM_eNVM_RW_0_ADDR[25] , 
        \eSRAM_eNVM_RW_0_ADDR[24] , \eSRAM_eNVM_RW_0_ADDR[23] , 
        \eSRAM_eNVM_RW_0_ADDR[22] , \eSRAM_eNVM_RW_0_ADDR[21] , 
        \eSRAM_eNVM_RW_0_ADDR[20] , \eSRAM_eNVM_RW_0_ADDR[19] , 
        \eSRAM_eNVM_RW_0_ADDR[18] , \eSRAM_eNVM_RW_0_ADDR[17] , 
        \eSRAM_eNVM_RW_0_ADDR[16] , \eSRAM_eNVM_RW_0_ADDR[15] , 
        \eSRAM_eNVM_RW_0_ADDR[14] , \eSRAM_eNVM_RW_0_ADDR[13] , 
        \eSRAM_eNVM_RW_0_ADDR[12] , \eSRAM_eNVM_RW_0_ADDR[11] , 
        \eSRAM_eNVM_RW_0_ADDR[10] , \eSRAM_eNVM_RW_0_ADDR[9] , 
        \eSRAM_eNVM_RW_0_ADDR[8] , \eSRAM_eNVM_RW_0_ADDR[7] , 
        \eSRAM_eNVM_RW_0_ADDR[6] , \eSRAM_eNVM_RW_0_ADDR[5] , 
        \eSRAM_eNVM_RW_0_ADDR[4] , \eSRAM_eNVM_RW_0_ADDR[3] , 
        \eSRAM_eNVM_RW_0_ADDR[2] }), .eSRAM_eNVM_access_0_FIC_0_CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .AHB_IF_0_VALID(AHB_IF_0_VALID), .AHB_IF_0_AHB_BUSY(
        AHB_IF_0_AHB_BUSY), .AHB_IF_0_BIF_1_HWRITE(
        AHB_IF_0_BIF_1_HWRITE), .HREADY_M_0_iv_i_0(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.HREADY_M_0_iv_i_0 )
        , .eSRAM_eNVM_RW_0_WRITE(eSRAM_eNVM_RW_0_WRITE), 
        .eSRAM_eNVM_RW_0_READ(eSRAM_eNVM_RW_0_READ), .N_546(N_546), 
        .defSlaveSMCurrentState(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMCurrentState )
        , .N_53(N_53), .defSlaveSMNextState(
        \eSRAM_eNVM_access_0.CoreAHBLite_0.matrix4x16.masterstage_0.default_slave_sm.defSlaveSMNextState )
        );
    OUTBUF \RD_obuf[7]  (.D(\RD_c[7] ), .PAD(RD[7]));
    OUTBUF \PRDATA_obuf[17]  (.D(\PRDATA_c[17] ), .PAD(PRDATA[17]));
    OUTBUF \PRDATA_obuf[3]  (.D(\PRDATA_c[3] ), .PAD(PRDATA[3]));
    OUTBUF \PRDATA_obuf[19]  (.D(\PRDATA_c[19] ), .PAD(PRDATA[19]));
    OUTBUF CS_obuf (.D(CS_c), .PAD(CS));
    OUTBUF \PRDATA_obuf[23]  (.D(\PRDATA_c[23] ), .PAD(PRDATA[23]));
    GND GND (.Y(GND_net_1));
    TRIBUFF CLKOUT_obuft (.D(CLKOUT_1), .E(CLKOUT_cl), .PAD(CLKOUT));
    OUTBUF \PRDATA_obuf[10]  (.D(\PRDATA_c[10] ), .PAD(PRDATA[10]));
    OUTBUF \PRDATA_obuf[12]  (.D(\PRDATA_c[12] ), .PAD(PRDATA[12]));
    OUTBUF \PRDATA_obuf[30]  (.D(\PRDATA_c[30] ), .PAD(PRDATA[30]));
    OUTBUF \PRDATA_obuf[16]  (.D(\PRDATA_c[16] ), .PAD(PRDATA[16]));
    OUTBUF \PRDATA_obuf[15]  (.D(\PRDATA_c[15] ), .PAD(PRDATA[15]));
    OUTBUF \PRDATA_obuf[0]  (.D(\PRDATA_c[0] ), .PAD(PRDATA[0]));
    OUTBUF \RD_obuf[0]  (.D(\RD_c[0] ), .PAD(RD[0]));
    OUTBUF \PRDATA_obuf[6]  (.D(\PRDATA_c[6] ), .PAD(PRDATA[6]));
    INBUF PWRITE_ibuf (.PAD(PWRITE), .Y(PWRITE_c));
    OUTBUF \PRDATA_obuf[5]  (.D(\PRDATA_c[5] ), .PAD(PRDATA[5]));
    OUTBUF \PRDATA_obuf[13]  (.D(\PRDATA_c[13] ), .PAD(PRDATA[13]));
    OUTBUF \PRDATA_obuf[9]  (.D(\PRDATA_c[9] ), .PAD(PRDATA[9]));
    OUTBUF \PRDATA_obuf[4]  (.D(\PRDATA_c[4] ), .PAD(PRDATA[4]));
    INBUF FAB_RESET_N_ibuf (.PAD(FAB_RESET_N), .Y(FAB_RESET_N_c));
    OUTBUF \RD_obuf[4]  (.D(\RD_c[4] ), .PAD(RD[4]));
    OUTBUF \RD_obuf[1]  (.D(\RD_c[1] ), .PAD(RD[1]));
    OUTBUF \PRDATA_obuf[24]  (.D(\PRDATA_c[24] ), .PAD(PRDATA[24]));
    OUTBUF \PRDATA_obuf[28]  (.D(\PRDATA_c[28] ), .PAD(PRDATA[28]));
    OUTBUF \RD_obuf[5]  (.D(\RD_c[5] ), .PAD(RD[5]));
    OUTBUF \PRDATA_obuf[7]  (.D(\PRDATA_c[7] ), .PAD(PRDATA[7]));
    SPI_Master SPI_Master_0 (.state({\SPI_Master_0.state[0] }), 
        .eSRAM_eNVM_RW_0_ram_waddr({\eSRAM_eNVM_RW_0_ram_waddr[4] , 
        \eSRAM_eNVM_RW_0_ram_waddr[3] , \eSRAM_eNVM_RW_0_ram_waddr[2] , 
        \eSRAM_eNVM_RW_0_ram_waddr[1] , \eSRAM_eNVM_RW_0_ram_waddr[0] })
        , .PRDATA_c({\PRDATA_c[31] , \PRDATA_c[30] , \PRDATA_c[29] , 
        \PRDATA_c[28] , \PRDATA_c[27] , \PRDATA_c[26] , \PRDATA_c[25] , 
        \PRDATA_c[24] , \PRDATA_c[23] , \PRDATA_c[22] , \PRDATA_c[21] , 
        \PRDATA_c[20] , \PRDATA_c[19] , \PRDATA_c[18] , \PRDATA_c[17] , 
        \PRDATA_c[16] , \PRDATA_c[15] , \PRDATA_c[14] , \PRDATA_c[13] , 
        \PRDATA_c[12] , \PRDATA_c[11] , \PRDATA_c[10] , \PRDATA_c[9] , 
        \PRDATA_c[8] , \PRDATA_c[7] , \PRDATA_c[6] , \PRDATA_c[5] , 
        \PRDATA_c[4] , \PRDATA_c[3] , \PRDATA_c[2] , \PRDATA_c[1] , 
        \PRDATA_c[0] }), .eSRAM_eNVM_RW_0_ram_wdata({
        \eSRAM_eNVM_RW_0_ram_wdata[31] , 
        \eSRAM_eNVM_RW_0_ram_wdata[30] , 
        \eSRAM_eNVM_RW_0_ram_wdata[29] , 
        \eSRAM_eNVM_RW_0_ram_wdata[28] , 
        \eSRAM_eNVM_RW_0_ram_wdata[27] , 
        \eSRAM_eNVM_RW_0_ram_wdata[26] , 
        \eSRAM_eNVM_RW_0_ram_wdata[25] , 
        \eSRAM_eNVM_RW_0_ram_wdata[24] , 
        \eSRAM_eNVM_RW_0_ram_wdata[23] , 
        \eSRAM_eNVM_RW_0_ram_wdata[22] , 
        \eSRAM_eNVM_RW_0_ram_wdata[21] , 
        \eSRAM_eNVM_RW_0_ram_wdata[20] , 
        \eSRAM_eNVM_RW_0_ram_wdata[19] , 
        \eSRAM_eNVM_RW_0_ram_wdata[18] , 
        \eSRAM_eNVM_RW_0_ram_wdata[17] , 
        \eSRAM_eNVM_RW_0_ram_wdata[16] , 
        \eSRAM_eNVM_RW_0_ram_wdata[15] , 
        \eSRAM_eNVM_RW_0_ram_wdata[14] , 
        \eSRAM_eNVM_RW_0_ram_wdata[13] , 
        \eSRAM_eNVM_RW_0_ram_wdata[12] , 
        \eSRAM_eNVM_RW_0_ram_wdata[11] , 
        \eSRAM_eNVM_RW_0_ram_wdata[10] , 
        \eSRAM_eNVM_RW_0_ram_wdata[9] , \eSRAM_eNVM_RW_0_ram_wdata[8] , 
        \eSRAM_eNVM_RW_0_ram_wdata[7] , \eSRAM_eNVM_RW_0_ram_wdata[6] , 
        \eSRAM_eNVM_RW_0_ram_wdata[5] , \eSRAM_eNVM_RW_0_ram_wdata[4] , 
        \eSRAM_eNVM_RW_0_ram_wdata[3] , \eSRAM_eNVM_RW_0_ram_wdata[2] , 
        \eSRAM_eNVM_RW_0_ram_wdata[1] , \eSRAM_eNVM_RW_0_ram_wdata[0] })
        , .PWRITE_c(PWRITE_c), .eSRAM_eNVM_access_0_FIC_0_CLK(
        eSRAM_eNVM_access_0_FIC_0_CLK), .MISO_c(MISO_c), 
        .eSRAM_eNVM_access_0_HPMS_READY(eSRAM_eNVM_access_0_HPMS_READY)
        , .CLKOUT_cl(CLKOUT_cl), .CLKOUT_1(CLKOUT_1), .MOSI_1(MOSI_1), 
        .ss_n_c(ss_n_c), .CS_c(CS_c), .MOSI_cl(MOSI_cl));
    OUTBUF \PRDATA_obuf[2]  (.D(\PRDATA_c[2] ), .PAD(PRDATA[2]));
    OUTBUF \PRDATA_obuf[21]  (.D(\PRDATA_c[21] ), .PAD(PRDATA[21]));
    
endmodule
